`default_nettype none
`include "fadd.sv"
/* verilator lint_off MULTITOP */
// hi
module fsqrt (input wire [31:0]  x,
             output wire [31:0] y,
             input clk);

    wire [31:0] a_table[1023:0];
    wire [31:0] b_table[1023:0];
    assign a_table = '{32'b00111110011101001111101000110010, 32'b00111110011101010001101101110101, 32'b00111110011101010011110011000110, 32'b00111110011101010101111000100100, 32'b00111110011101010111111110001111, 32'b00111110011101011010000100001001, 32'b00111110011101011100001010010000, 32'b00111110011101011110010000100101, 32'b00111110011101100000010111000111, 32'b00111110011101100010011101111000, 32'b00111110011101100100100100110110, 32'b00111110011101100110101100000010, 32'b00111110011101101000110011011100, 32'b00111110011101101010111011000100, 32'b00111110011101101101000010111010, 32'b00111110011101101111001010111110, 32'b00111110011101110001010011010001, 32'b00111110011101110011011011110001, 32'b00111110011101110101100100011111, 32'b00111110011101110111101101011100, 32'b00111110011101111001110110100111, 32'b00111110011101111100000000000000, 32'b00111110011101111110001001101000, 32'b00111110011110000000010011011101, 32'b00111110011110000010011101100010, 32'b00111110011110000100100111110100, 32'b00111110011110000110110010010101, 32'b00111110011110001000111101000101, 32'b00111110011110001011001000000011, 32'b00111110011110001101010011010000, 32'b00111110011110001111011110101011, 32'b00111110011110010001101010010101, 32'b00111110011110010011110110001110, 32'b00111110011110010110000010010101, 32'b00111110011110011000001110101011, 32'b00111110011110011010011011010001, 32'b00111110011110011100101000000100, 32'b00111110011110011110110101000111, 32'b00111110011110100001000010011001, 32'b00111110011110100011001111111010, 32'b00111110011110100101011101101010, 32'b00111110011110100111101011101001, 32'b00111110011110101001111001110111, 32'b00111110011110101100001000010100, 32'b00111110011110101110010111000000, 32'b00111110011110110000100101111100, 32'b00111110011110110010110101000111, 32'b00111110011110110101000100100001, 32'b00111110011110110111010100001010, 32'b00111110011110111001100100000011, 32'b00111110011110111011110100001100, 32'b00111110011110111110000100100100, 32'b00111110011111000000010101001011, 32'b00111110011111000010100110000010, 32'b00111110011111000100110111001001, 32'b00111110011111000111001000011111, 32'b00111110011111001001011010000110, 32'b00111110011111001011101011111011, 32'b00111110011111001101111110000001, 32'b00111110011111010000010000010111, 32'b00111110011111010010100010111100, 32'b00111110011111010100110101110001, 32'b00111110011111010111001000110111, 32'b00111110011111011001011100001100, 32'b00111110011111011011101111110010, 32'b00111110011111011110000011100111, 32'b00111110011111100000010111101101, 32'b00111110011111100010101100000011, 32'b00111110011111100101000000101001, 32'b00111110011111100111010101100000, 32'b00111110011111101001101010100111, 32'b00111110011111101011111111111110, 32'b00111110011111101110010101100110, 32'b00111110011111110000101011011110, 32'b00111110011111110011000001100111, 32'b00111110011111110101011000000000, 32'b00111110011111110111101110101010, 32'b00111110011111111010000101100101, 32'b00111110011111111100011100110000, 32'b00111110011111111110110100001100, 32'b00111110100000000000100101111101, 32'b00111110100000000001110001111100, 32'b00111110100000000010111110000011, 32'b00111110100000000100001010010011, 32'b00111110100000000101010110101011, 32'b00111110100000000110100011001100, 32'b00111110100000000111101111110110, 32'b00111110100000001000111100101000, 32'b00111110100000001010001001100011, 32'b00111110100000001011010110100110, 32'b00111110100000001100100011110010, 32'b00111110100000001101110001000111, 32'b00111110100000001110111110100100, 32'b00111110100000010000001100001011, 32'b00111110100000010001011001111001, 32'b00111110100000010010100111110001, 32'b00111110100000010011110101110010, 32'b00111110100000010101000011111011, 32'b00111110100000010110010010001101, 32'b00111110100000010111100000101001, 32'b00111110100000011000101111001101, 32'b00111110100000011001111101111010, 32'b00111110100000011011001100110000, 32'b00111110100000011100011011101111, 32'b00111110100000011101101010110111, 32'b00111110100000011110111010001000, 32'b00111110100000100000001001100010, 32'b00111110100000100001011001000101, 32'b00111110100000100010101000110010, 32'b00111110100000100011111000100111, 32'b00111110100000100101001000100110, 32'b00111110100000100110011000101110, 32'b00111110100000100111101001000000, 32'b00111110100000101000111001011010, 32'b00111110100000101010001001111110, 32'b00111110100000101011011010101011, 32'b00111110100000101100101011100010, 32'b00111110100000101101111100100010, 32'b00111110100000101111001101101011, 32'b00111110100000110000011110111110, 32'b00111110100000110001110000011010, 32'b00111110100000110011000010000000, 32'b00111110100000110100010011101111, 32'b00111110100000110101100101101000, 32'b00111110100000110110110111101010, 32'b00111110100000111000001001110110, 32'b00111110100000111001011100001100, 32'b00111110100000111010101110101011, 32'b00111110100000111100000001010101, 32'b00111110100000111101010100000111, 32'b00111110100000111110100111000100, 32'b00111110100000111111111010001010, 32'b00111110100001000001001101011011, 32'b00111110100001000010100000110101, 32'b00111110100001000011110100011001, 32'b00111110100001000101001000000111, 32'b00111110100001000110011011111110, 32'b00111110100001000111110000000000, 32'b00111110100001001001000100001100, 32'b00111110100001001010011000100010, 32'b00111110100001001011101101000010, 32'b00111110100001001101000001101100, 32'b00111110100001001110010110100000, 32'b00111110100001001111101011011111, 32'b00111110100001010001000000100111, 32'b00111110100001010010010101111010, 32'b00111110100001010011101011010111, 32'b00111110100001010101000000111110, 32'b00111110100001010110010110110000, 32'b00111110100001010111101100101100, 32'b00111110100001011001000010110011, 32'b00111110100001011010011001000011, 32'b00111110100001011011101111011111, 32'b00111110100001011101000110000101, 32'b00111110100001011110011100110101, 32'b00111110100001011111110011110000, 32'b00111110100001100001001010110101, 32'b00111110100001100010100010000101, 32'b00111110100001100011111001100000, 32'b00111110100001100101010001000110, 32'b00111110100001100110101000110110, 32'b00111110100001101000000000110001, 32'b00111110100001101001011000110111, 32'b00111110100001101010110001000111, 32'b00111110100001101100001001100011, 32'b00111110100001101101100010001001, 32'b00111110100001101110111010111010, 32'b00111110100001110000010011110111, 32'b00111110100001110001101100111110, 32'b00111110100001110011000110010000, 32'b00111110100001110100011111101110, 32'b00111110100001110101111001010110, 32'b00111110100001110111010011001010, 32'b00111110100001111000101101001001, 32'b00111110100001111010000111010011, 32'b00111110100001111011100001101000, 32'b00111110100001111100111100001001, 32'b00111110100001111110010110110101, 32'b00111110100001111111110001101100, 32'b00111110100010000001001100101111, 32'b00111110100010000010100111111101, 32'b00111110100010000100000011010110, 32'b00111110100010000101011110111100, 32'b00111110100010000110111010101100, 32'b00111110100010001000010110101001, 32'b00111110100010001001110010110001, 32'b00111110100010001011001111000100, 32'b00111110100010001100101011100100, 32'b00111110100010001110001000001111, 32'b00111110100010001111100101000110, 32'b00111110100010010001000010001000, 32'b00111110100010010010011111010111, 32'b00111110100010010011111100110001, 32'b00111110100010010101011010011000, 32'b00111110100010010110111000001010, 32'b00111110100010011000010110001001, 32'b00111110100010011001110100010011, 32'b00111110100010011011010010101010, 32'b00111110100010011100110001001100, 32'b00111110100010011110001111111011, 32'b00111110100010011111101110110110, 32'b00111110100010100001001101111110, 32'b00111110100010100010101101010010, 32'b00111110100010100100001100110010, 32'b00111110100010100101101100011110, 32'b00111110100010100111001100010111, 32'b00111110100010101000101100011101, 32'b00111110100010101010001100101110, 32'b00111110100010101011101101001101, 32'b00111110100010101101001101111000, 32'b00111110100010101110101110110000, 32'b00111110100010110000001111110100, 32'b00111110100010110001110001000101, 32'b00111110100010110011010010100011, 32'b00111110100010110100110100001110, 32'b00111110100010110110010110000110, 32'b00111110100010110111111000001010, 32'b00111110100010111001011010011100, 32'b00111110100010111010111100111010, 32'b00111110100010111100011111100110, 32'b00111110100010111110000010011110, 32'b00111110100010111111100101100100, 32'b00111110100011000001001000110111, 32'b00111110100011000010101100010111, 32'b00111110100011000100010000000101, 32'b00111110100011000101110011111111, 32'b00111110100011000111011000000111, 32'b00111110100011001000111100011101, 32'b00111110100011001010100001000000, 32'b00111110100011001100000101110000, 32'b00111110100011001101101010101110, 32'b00111110100011001111001111111010, 32'b00111110100011010000110101010011, 32'b00111110100011010010011010111010, 32'b00111110100011010100000000101111, 32'b00111110100011010101100110110010, 32'b00111110100011010111001101000010, 32'b00111110100011011000110011100000, 32'b00111110100011011010011010001100, 32'b00111110100011011100000001000111, 32'b00111110100011011101101000001111, 32'b00111110100011011111001111100101, 32'b00111110100011100000110111001010, 32'b00111110100011100010011110111100, 32'b00111110100011100100000110111101, 32'b00111110100011100101101111001100, 32'b00111110100011100111010111101010, 32'b00111110100011101001000000010110, 32'b00111110100011101010101001010000, 32'b00111110100011101100010010011001, 32'b00111110100011101101111011110000, 32'b00111110100011101111100101010110, 32'b00111110100011110001001111001011, 32'b00111110100011110010111001001110, 32'b00111110100011110100100011100000, 32'b00111110100011110110001110000001, 32'b00111110100011110111111000110001, 32'b00111110100011111001100011110000, 32'b00111110100011111011001110111101, 32'b00111110100011111100111010011010, 32'b00111110100011111110100110000110, 32'b00111110100100000000010010000001, 32'b00111110100100000001111110001011, 32'b00111110100100000011101010100100, 32'b00111110100100000101010111001101, 32'b00111110100100000111000100000101, 32'b00111110100100001000110001001101, 32'b00111110100100001010011110100100, 32'b00111110100100001100001100001010, 32'b00111110100100001101111010000000, 32'b00111110100100001111101000000110, 32'b00111110100100010001010110011011, 32'b00111110100100010011000101000001, 32'b00111110100100010100110011110110, 32'b00111110100100010110100010111011, 32'b00111110100100011000010010010000, 32'b00111110100100011010000001110100, 32'b00111110100100011011110001101001, 32'b00111110100100011101100001101110, 32'b00111110100100011111010010000100, 32'b00111110100100100001000010101001, 32'b00111110100100100010110011011111, 32'b00111110100100100100100100100101, 32'b00111110100100100110010101111100, 32'b00111110100100101000000111100011, 32'b00111110100100101001111001011011, 32'b00111110100100101011101011100011, 32'b00111110100100101101011101111100, 32'b00111110100100101111010000100110, 32'b00111110100100110001000011100000, 32'b00111110100100110010110110101100, 32'b00111110100100110100101010001000, 32'b00111110100100110110011101110101, 32'b00111110100100111000010001110100, 32'b00111110100100111010000110000011, 32'b00111110100100111011111010100100, 32'b00111110100100111101101111010110, 32'b00111110100100111111100100011001, 32'b00111110100101000001011001101110, 32'b00111110100101000011001111010100, 32'b00111110100101000101000101001100, 32'b00111110100101000110111011010110, 32'b00111110100101001000110001110001, 32'b00111110100101001010101000011101, 32'b00111110100101001100011111011100, 32'b00111110100101001110010110101100, 32'b00111110100101010000001110001111, 32'b00111110100101010010000110000011, 32'b00111110100101010011111110001010, 32'b00111110100101010101110110100011, 32'b00111110100101010111101111001110, 32'b00111110100101011001101000001011, 32'b00111110100101011011100001011010, 32'b00111110100101011101011010111101, 32'b00111110100101011111010100110001, 32'b00111110100101100001001110111000, 32'b00111110100101100011001001010010, 32'b00111110100101100101000011111111, 32'b00111110100101100110111110111110, 32'b00111110100101101000111010010001, 32'b00111110100101101010110101110110, 32'b00111110100101101100110001101111, 32'b00111110100101101110101101111010, 32'b00111110100101110000101010011001, 32'b00111110100101110010100111001011, 32'b00111110100101110100100100010000, 32'b00111110100101110110100001101001, 32'b00111110100101111000011111010101, 32'b00111110100101111010011101010101, 32'b00111110100101111100011011101001, 32'b00111110100101111110011010010000, 32'b00111110100110000000011001001011, 32'b00111110100110000010011000011010, 32'b00111110100110000100010111111110, 32'b00111110100110000110010111110101, 32'b00111110100110001000011000000000, 32'b00111110100110001010011000100000, 32'b00111110100110001100011001010100, 32'b00111110100110001110011010011100, 32'b00111110100110010000011011111001, 32'b00111110100110010010011101101010, 32'b00111110100110010100011111110000, 32'b00111110100110010110100010001011, 32'b00111110100110011000100100111011, 32'b00111110100110011010100111111111, 32'b00111110100110011100101011011001, 32'b00111110100110011110101111001000, 32'b00111110100110100000110011001100, 32'b00111110100110100010110111100101, 32'b00111110100110100100111100010011, 32'b00111110100110100111000001011000, 32'b00111110100110101001000110110001, 32'b00111110100110101011001100100000, 32'b00111110100110101101010010100101, 32'b00111110100110101111011001000000, 32'b00111110100110110001011111110001, 32'b00111110100110110011100110110111, 32'b00111110100110110101101110010100, 32'b00111110100110110111110110000111, 32'b00111110100110111001111110010001, 32'b00111110100110111100000110110000, 32'b00111110100110111110001111100111, 32'b00111110100111000000011000110011, 32'b00111110100111000010100010010111, 32'b00111110100111000100101100010001, 32'b00111110100111000110110110100010, 32'b00111110100111001001000001001010, 32'b00111110100111001011001100001001, 32'b00111110100111001101010111100000, 32'b00111110100111001111100011001101, 32'b00111110100111010001101111010010, 32'b00111110100111010011111011101111, 32'b00111110100111010110001000100011, 32'b00111110100111011000010101101110, 32'b00111110100111011010100011010010, 32'b00111110100111011100110001001101, 32'b00111110100111011110111111100001, 32'b00111110100111100001001110001100, 32'b00111110100111100011011101010000, 32'b00111110100111100101101100101100, 32'b00111110100111100111111100100001, 32'b00111110100111101010001100101110, 32'b00111110100111101100011101010011, 32'b00111110100111101110101110010010, 32'b00111110100111110000111111101001, 32'b00111110100111110011010001011001, 32'b00111110100111110101100011100010, 32'b00111110100111110111110110000101, 32'b00111110100111111010001001000001, 32'b00111110100111111100011100010110, 32'b00111110100111111110110000000101, 32'b00111110101000000001000100001101, 32'b00111110101000000011011000110000, 32'b00111110101000000101101101101100, 32'b00111110101000001000000011000010, 32'b00111110101000001010011000110010, 32'b00111110101000001100101110111101, 32'b00111110101000001111000101100001, 32'b00111110101000010001011100100001, 32'b00111110101000010011110011111011, 32'b00111110101000010110001011101111, 32'b00111110101000011000100011111111, 32'b00111110101000011010111100101010, 32'b00111110101000011101010101101111, 32'b00111110101000011111101111010000, 32'b00111110101000100010001001001100, 32'b00111110101000100100100011100100, 32'b00111110101000100110111110010111, 32'b00111110101000101001011001100110, 32'b00111110101000101011110101010001, 32'b00111110101000101110010001011000, 32'b00111110101000110000101101111011, 32'b00111110101000110011001010111011, 32'b00111110101000110101101000010110, 32'b00111110101000111000000110001110, 32'b00111110101000111010100100100011, 32'b00111110101000111101000011010101, 32'b00111110101000111111100010100100, 32'b00111110101001000010000010001111, 32'b00111110101001000100100010011000, 32'b00111110101001000111000010111111, 32'b00111110101001001001100100000010, 32'b00111110101001001100000101100100, 32'b00111110101001001110100111100011, 32'b00111110101001010001001010000000, 32'b00111110101001010011101100111011, 32'b00111110101001010110010000010101, 32'b00111110101001011000110100001100, 32'b00111110101001011011011000100011, 32'b00111110101001011101111101010111, 32'b00111110101001100000100010101011, 32'b00111110101001100011001000011110, 32'b00111110101001100101101110110000, 32'b00111110101001101000010101100000, 32'b00111110101001101010111100110001, 32'b00111110101001101101100100100001, 32'b00111110101001110000001100110001, 32'b00111110101001110010110101100000, 32'b00111110101001110101011110110000, 32'b00111110101001111000001000011111, 32'b00111110101001111010110010101111, 32'b00111110101001111101011101100000, 32'b00111110101010000000001000110001, 32'b00111110101010000010110100100100, 32'b00111110101010000101100000110111, 32'b00111110101010001000001101101011, 32'b00111110101010001010111011000001, 32'b00111110101010001101101000111000, 32'b00111110101010010000010111010000, 32'b00111110101010010011000110001011, 32'b00111110101010010101110101101000, 32'b00111110101010011000100101100111, 32'b00111110101010011011010110001000, 32'b00111110101010011110000111001011, 32'b00111110101010100000111000110010, 32'b00111110101010100011101010111011, 32'b00111110101010100110011101100111, 32'b00111110101010101001010000110111, 32'b00111110101010101100000100101010, 32'b00111110101010101110111001000001, 32'b00111110101010110001101101111011, 32'b00111110101010110100100011011010, 32'b00111110101010110111011001011100, 32'b00111110101010111010010000000011, 32'b00111110101010111101000111001110, 32'b00111110101010111111111110111111, 32'b00111110101011000010110111010100, 32'b00111110101011000101110000001110, 32'b00111110101011001000101001101110, 32'b00111110101011001011100011110011, 32'b00111110101011001110011110011101, 32'b00111110101011010001011001101110, 32'b00111110101011010100010101100101, 32'b00111110101011010111010010000010, 32'b00111110101011011010001111000101, 32'b00111110101011011101001100110000, 32'b00111110101011100000001011000001, 32'b00111110101011100011001001111001, 32'b00111110101011100110001001011001, 32'b00111110101011101001001001100000, 32'b00111110101011101100001010001111, 32'b00111110101011101111001011100110, 32'b00111110101011110010001101100110, 32'b00111110101011110101010000001101, 32'b00111110101011111000010011011101, 32'b00111110101011111011010111010111, 32'b00111110101011111110011011111001, 32'b00111110101100000001100001000100, 32'b00111110101100000100100110111001, 32'b00111110101100000111101101011000, 32'b00111110101100001010110100100001, 32'b00111110101100001101111100010100, 32'b00111110101100010001000100110010, 32'b00111110101100010100001101111010, 32'b00111110101100010111010111101101, 32'b00111110101100011010100010001011, 32'b00111110101100011101101101010101, 32'b00111110101100100000111001001010, 32'b00111110101100100100000101101100, 32'b00111110101100100111010010111001, 32'b00111110101100101010100000110011, 32'b00111110101100101101101111011001, 32'b00111110101100110000111110101101, 32'b00111110101100110100001110101101, 32'b00111110101100110111011111011011, 32'b00111110101100111010110000110111, 32'b00111110101100111110000011000000, 32'b00111110101101000001010101111000, 32'b00111110101101000100101001011110, 32'b00111110101101000111111101110011, 32'b00111110101101001011010010110111, 32'b00111110101101001110101000101010, 32'b00111110101101010001000001000101, 32'b00111110101101010010011011101110, 32'b00111110101101010011110110100000, 32'b00111110101101010101010001011010, 32'b00111110101101010110101100011101, 32'b00111110101101011000000111101000, 32'b00111110101101011001100010111100, 32'b00111110101101011010111110011000, 32'b00111110101101011100011001111101, 32'b00111110101101011101110101101011, 32'b00111110101101011111010001100010, 32'b00111110101101100000101101100001, 32'b00111110101101100010001001101001, 32'b00111110101101100011100101111010, 32'b00111110101101100101000010010011, 32'b00111110101101100110011110110101, 32'b00111110101101100111111011100001, 32'b00111110101101101001011000010100, 32'b00111110101101101010110101010001, 32'b00111110101101101100010010010111, 32'b00111110101101101101101111100110, 32'b00111110101101101111001100111101, 32'b00111110101101110000101010011101, 32'b00111110101101110010001000000111, 32'b00111110101101110011100101111001, 32'b00111110101101110101000011110101, 32'b00111110101101110110100001111001, 32'b00111110101101111000000000000111, 32'b00111110101101111001011110011101, 32'b00111110101101111010111100111101, 32'b00111110101101111100011011100110, 32'b00111110101101111101111010011000, 32'b00111110101101111111011001010011, 32'b00111110101110000000111000010111, 32'b00111110101110000010010111100101, 32'b00111110101110000011110110111100, 32'b00111110101110000101010110011100, 32'b00111110101110000110110110000101, 32'b00111110101110001000010101111000, 32'b00111110101110001001110101110100, 32'b00111110101110001011010101111001, 32'b00111110101110001100110110001000, 32'b00111110101110001110010110100000, 32'b00111110101110001111110111000010, 32'b00111110101110010001010111101101, 32'b00111110101110010010111000100001, 32'b00111110101110010100011001100000, 32'b00111110101110010101111010100111, 32'b00111110101110010111011011111000, 32'b00111110101110011000111101010011, 32'b00111110101110011010011110110111, 32'b00111110101110011100000000100101, 32'b00111110101110011101100010011101, 32'b00111110101110011111000100011110, 32'b00111110101110100000100110101001, 32'b00111110101110100010001000111110, 32'b00111110101110100011101011011101, 32'b00111110101110100101001110000101, 32'b00111110101110100110110000110111, 32'b00111110101110101000010011110011, 32'b00111110101110101001110110111001, 32'b00111110101110101011011010001000, 32'b00111110101110101100111101100010, 32'b00111110101110101110100001000101, 32'b00111110101110110000000100110011, 32'b00111110101110110001101000101010, 32'b00111110101110110011001100101011, 32'b00111110101110110100110000110111, 32'b00111110101110110110010101001100, 32'b00111110101110110111111001101100, 32'b00111110101110111001011110010110, 32'b00111110101110111011000011001010, 32'b00111110101110111100101000001000, 32'b00111110101110111110001101010000, 32'b00111110101110111111110010100010, 32'b00111110101111000001010111111111, 32'b00111110101111000010111101100110, 32'b00111110101111000100100011010111, 32'b00111110101111000110001001010011, 32'b00111110101111000111101111011001, 32'b00111110101111001001010101101001, 32'b00111110101111001010111100000100, 32'b00111110101111001100100010101001, 32'b00111110101111001110001001011001, 32'b00111110101111001111110000010011, 32'b00111110101111010001010111011000, 32'b00111110101111010010111110100111, 32'b00111110101111010100100110000001, 32'b00111110101111010110001101100101, 32'b00111110101111010111110101010100, 32'b00111110101111011001011101001110, 32'b00111110101111011011000101010011, 32'b00111110101111011100101101100010, 32'b00111110101111011110010101111100, 32'b00111110101111011111111110100000, 32'b00111110101111100001100111010000, 32'b00111110101111100011010000001010, 32'b00111110101111100100111001001111, 32'b00111110101111100110100010011111, 32'b00111110101111101000001011111011, 32'b00111110101111101001110101100000, 32'b00111110101111101011011111010001, 32'b00111110101111101101001001001101, 32'b00111110101111101110110011010100, 32'b00111110101111110000011101100111, 32'b00111110101111110010001000000100, 32'b00111110101111110011110010101100, 32'b00111110101111110101011101100000, 32'b00111110101111110111001000011110, 32'b00111110101111111000110011101000, 32'b00111110101111111010011110111101, 32'b00111110101111111100001010011110, 32'b00111110101111111101110110001010, 32'b00111110101111111111100010000001, 32'b00111110110000000001001110000011, 32'b00111110110000000010111010010001, 32'b00111110110000000100100110101011, 32'b00111110110000000110010011010000, 32'b00111110110000001000000000000000, 32'b00111110110000001001101100111100, 32'b00111110110000001011011010000011, 32'b00111110110000001101000111010111, 32'b00111110110000001110110100110101, 32'b00111110110000010000100010100000, 32'b00111110110000010010010000010110, 32'b00111110110000010011111110011000, 32'b00111110110000010101101100100101, 32'b00111110110000010111011010111111, 32'b00111110110000011001001001100100, 32'b00111110110000011010111000010101, 32'b00111110110000011100100111010010, 32'b00111110110000011110010110011011, 32'b00111110110000100000000101110000, 32'b00111110110000100001110101010001, 32'b00111110110000100011100100111101, 32'b00111110110000100101010100110110, 32'b00111110110000100111000100111100, 32'b00111110110000101000110101001101, 32'b00111110110000101010100101101010, 32'b00111110110000101100010110010100, 32'b00111110110000101110000111001010, 32'b00111110110000101111111000001100, 32'b00111110110000110001101001011010, 32'b00111110110000110011011010110101, 32'b00111110110000110101001100011100, 32'b00111110110000110110111110001111, 32'b00111110110000111000110000001111, 32'b00111110110000111010100010011100, 32'b00111110110000111100010100110101, 32'b00111110110000111110000111011010, 32'b00111110110000111111111010001100, 32'b00111110110001000001101101001011, 32'b00111110110001000011100000010111, 32'b00111110110001000101010011101111, 32'b00111110110001000111000111010100, 32'b00111110110001001000111011000101, 32'b00111110110001001010101111000100, 32'b00111110110001001100100011001111, 32'b00111110110001001110010111100111, 32'b00111110110001010000001100001100, 32'b00111110110001010010000000111110, 32'b00111110110001010011110101111101, 32'b00111110110001010101101011001001, 32'b00111110110001010111100000100010, 32'b00111110110001011001010110001000, 32'b00111110110001011011001011111100, 32'b00111110110001011101000001111100, 32'b00111110110001011110111000001010, 32'b00111110110001100000101110100101, 32'b00111110110001100010100101001110, 32'b00111110110001100100011100000011, 32'b00111110110001100110010011000110, 32'b00111110110001101000001010010111, 32'b00111110110001101010000001110101, 32'b00111110110001101011111001100000, 32'b00111110110001101101110001011001, 32'b00111110110001101111101001100000, 32'b00111110110001110001100001110100, 32'b00111110110001110011011010010110, 32'b00111110110001110101010011000101, 32'b00111110110001110111001100000010, 32'b00111110110001111001000101001101, 32'b00111110110001111010111110100110, 32'b00111110110001111100111000001101, 32'b00111110110001111110110010000010, 32'b00111110110010000000101100000100, 32'b00111110110010000010100110010101, 32'b00111110110010000100100000110011, 32'b00111110110010000110011011100000, 32'b00111110110010001000010110011011, 32'b00111110110010001010010001100100, 32'b00111110110010001100001100111011, 32'b00111110110010001110001000100000, 32'b00111110110010010000000100010100, 32'b00111110110010010010000000010110, 32'b00111110110010010011111100100110, 32'b00111110110010010101111001000101, 32'b00111110110010010111110101110010, 32'b00111110110010011001110010101110, 32'b00111110110010011011101111111000, 32'b00111110110010011101101101010001, 32'b00111110110010011111101010111000, 32'b00111110110010100001101000101110, 32'b00111110110010100011100110110011, 32'b00111110110010100101100101000110, 32'b00111110110010100111100011101001, 32'b00111110110010101001100010011010, 32'b00111110110010101011100001011010, 32'b00111110110010101101100000101001, 32'b00111110110010101111100000000111, 32'b00111110110010110001011111110101, 32'b00111110110010110011011111110001, 32'b00111110110010110101011111111100, 32'b00111110110010110111100000010111, 32'b00111110110010111001100001000000, 32'b00111110110010111011100001111001, 32'b00111110110010111101100011000010, 32'b00111110110010111111100100011010, 32'b00111110110011000001100110000001, 32'b00111110110011000011100111110111, 32'b00111110110011000101101001111101, 32'b00111110110011000111101100010011, 32'b00111110110011001001101110111000, 32'b00111110110011001011110001101101, 32'b00111110110011001101110100110010, 32'b00111110110011001111111000000110, 32'b00111110110011010001111011101010, 32'b00111110110011010011111111011110, 32'b00111110110011010110000011100010, 32'b00111110110011011000000111110110, 32'b00111110110011011010001100011010, 32'b00111110110011011100010001001110, 32'b00111110110011011110010110010010, 32'b00111110110011100000011011100110, 32'b00111110110011100010100001001010, 32'b00111110110011100100100110111111, 32'b00111110110011100110101101000100, 32'b00111110110011101000110011011001, 32'b00111110110011101010111001111111, 32'b00111110110011101101000000110101, 32'b00111110110011101111000111111100, 32'b00111110110011110001001111010011, 32'b00111110110011110011010110111011, 32'b00111110110011110101011110110100, 32'b00111110110011110111100110111101, 32'b00111110110011111001101111010111, 32'b00111110110011111011111000000010, 32'b00111110110011111110000000111110, 32'b00111110110100000000001010001011, 32'b00111110110100000010010011101001, 32'b00111110110100000100011101010111, 32'b00111110110100000110100111010111, 32'b00111110110100001000110001101000, 32'b00111110110100001010111100001011, 32'b00111110110100001101000110111110, 32'b00111110110100001111010010000011, 32'b00111110110100010001011101011010, 32'b00111110110100010011101001000001, 32'b00111110110100010101110100111011, 32'b00111110110100011000000001000101, 32'b00111110110100011010001101100010, 32'b00111110110100011100011010010000, 32'b00111110110100011110100111010000, 32'b00111110110100100000110100100010, 32'b00111110110100100011000010000101, 32'b00111110110100100101001111111010, 32'b00111110110100100111011110000010, 32'b00111110110100101001101100011011, 32'b00111110110100101011111011000111, 32'b00111110110100101110001010000100, 32'b00111110110100110000011001010100, 32'b00111110110100110010101000110110, 32'b00111110110100110100111000101011, 32'b00111110110100110111001000110010, 32'b00111110110100111001011001001011, 32'b00111110110100111011101001110111, 32'b00111110110100111101111010110101, 32'b00111110110101000000001100000110, 32'b00111110110101000010011101101010, 32'b00111110110101000100101111100001, 32'b00111110110101000111000001101010, 32'b00111110110101001001010100000110, 32'b00111110110101001011100110110101, 32'b00111110110101001101111001110111, 32'b00111110110101010000001101001101, 32'b00111110110101010010100000110101, 32'b00111110110101010100110100110001, 32'b00111110110101010111001001000000, 32'b00111110110101011001011101100010, 32'b00111110110101011011110010010111, 32'b00111110110101011110000111100001, 32'b00111110110101100000011100111101, 32'b00111110110101100010110010101101, 32'b00111110110101100101001000110001, 32'b00111110110101100111011111001001, 32'b00111110110101101001110101110101, 32'b00111110110101101100001100110100, 32'b00111110110101101110100100000111, 32'b00111110110101110000111011101111, 32'b00111110110101110011010011101010, 32'b00111110110101110101101011111001, 32'b00111110110101111000000100011101, 32'b00111110110101111010011101010101, 32'b00111110110101111100110110100010, 32'b00111110110101111111010000000011, 32'b00111110110110000001101001111000, 32'b00111110110110000100000100000010, 32'b00111110110110000110011110100000, 32'b00111110110110001000111001010100, 32'b00111110110110001011010100011100, 32'b00111110110110001101101111111001, 32'b00111110110110010000001011101011, 32'b00111110110110010010100111110010, 32'b00111110110110010101000100001110, 32'b00111110110110010111100000111111, 32'b00111110110110011001111110000101, 32'b00111110110110011100011011100001, 32'b00111110110110011110111001010010, 32'b00111110110110100001010111011001, 32'b00111110110110100011110101110101, 32'b00111110110110100110010100100110, 32'b00111110110110101000110011101110, 32'b00111110110110101011010011001011, 32'b00111110110110101101110010111110, 32'b00111110110110110000010011000111, 32'b00111110110110110010110011100110, 32'b00111110110110110101010100011011, 32'b00111110110110110111110101100110, 32'b00111110110110111010010111000111, 32'b00111110110110111100111000111111, 32'b00111110110110111111011011001101, 32'b00111110110111000001111101110010, 32'b00111110110111000100100000101101, 32'b00111110110111000111000011111111, 32'b00111110110111001001100111100111, 32'b00111110110111001100001011100111, 32'b00111110110111001110101111111101, 32'b00111110110111010001010100101010, 32'b00111110110111010011111001101110, 32'b00111110110111010110011111001010, 32'b00111110110111011001000100111100, 32'b00111110110111011011101011000110, 32'b00111110110111011110010001101000, 32'b00111110110111100000111000100000, 32'b00111110110111100011011111110001, 32'b00111110110111100110000111011001, 32'b00111110110111101000101111011001, 32'b00111110110111101011010111110000, 32'b00111110110111101110000000100000, 32'b00111110110111110000101001100111, 32'b00111110110111110011010011000111, 32'b00111110110111110101111100111111, 32'b00111110110111111000100111001111, 32'b00111110110111111011010001110111, 32'b00111110110111111101111100111000, 32'b00111110111000000000101000010010, 32'b00111110111000000011010100000100, 32'b00111110111000000110000000001111, 32'b00111110111000001000101100110010, 32'b00111110111000001011011001101111, 32'b00111110111000001110000111000101, 32'b00111110111000010000110100110011, 32'b00111110111000010011100010111011, 32'b00111110111000010110010001011100, 32'b00111110111000011001000000010111, 32'b00111110111000011011101111101011, 32'b00111110111000011110011111011001, 32'b00111110111000100001001111100000, 32'b00111110111000100100000000000001, 32'b00111110111000100110110000111100, 32'b00111110111000101001100010010001, 32'b00111110111000101100010100000001, 32'b00111110111000101111000110001010, 32'b00111110111000110001111000101101, 32'b00111110111000110100101011101011, 32'b00111110111000110111011111000100, 32'b00111110111000111010010010110111, 32'b00111110111000111101000111000101, 32'b00111110111000111111111011101101, 32'b00111110111001000010110000110000, 32'b00111110111001000101100110001111, 32'b00111110111001001000011100001000, 32'b00111110111001001011010010011101, 32'b00111110111001001110001001001101, 32'b00111110111001010001000000011000, 32'b00111110111001010011110111111111, 32'b00111110111001010110110000000010, 32'b00111110111001011001101000100000, 32'b00111110111001011100100001011011, 32'b00111110111001011111011010110001, 32'b00111110111001100010010100100011, 32'b00111110111001100101001110110010, 32'b00111110111001101000001001011100, 32'b00111110111001101011000100100011, 32'b00111110111001101110000000000111, 32'b00111110111001110000111100000111, 32'b00111110111001110011111000100101, 32'b00111110111001110110110101011110, 32'b00111110111001111001110010110101, 32'b00111110111001111100110000101001, 32'b00111110111001111111101110111011, 32'b00111110111010000010101101101001, 32'b00111110111010000101101100110101, 32'b00111110111010001000101100011111, 32'b00111110111010001011101100100110, 32'b00111110111010001110101101001011, 32'b00111110111010010001101110001110, 32'b00111110111010010100101111101111, 32'b00111110111010010111110001101110, 32'b00111110111010011010110100001100, 32'b00111110111010011101110111001000, 32'b00111110111010100000111010100010, 32'b00111110111010100011111110011011, 32'b00111110111010100111000010110011, 32'b00111110111010101010000111101010, 32'b00111110111010101101001101000000, 32'b00111110111010110000010010110101, 32'b00111110111010110011011001001001, 32'b00111110111010110110011111111101, 32'b00111110111010111001100111010001, 32'b00111110111010111100101111000100, 32'b00111110111010111111110111010110, 32'b00111110111011000011000000001001, 32'b00111110111011000110001001011100, 32'b00111110111011001001010011001111, 32'b00111110111011001100011101100011, 32'b00111110111011001111101000010111, 32'b00111110111011010010110011101011, 32'b00111110111011010101111111100001, 32'b00111110111011011001001011110111, 32'b00111110111011011100011000101110, 32'b00111110111011011111100110000111, 32'b00111110111011100010110100000000, 32'b00111110111011100110000010011100, 32'b00111110111011101001010001011001, 32'b00111110111011101100100000110111, 32'b00111110111011101111110000111000, 32'b00111110111011110011000001011010, 32'b00111110111011110110010010011111, 32'b00111110111011111001100100000110, 32'b00111110111011111100110110001111, 32'b00111110111100000000001000111011, 32'b00111110111100000011011100001010, 32'b00111110111100000110101111111100, 32'b00111110111100001010000100010001, 32'b00111110111100001101011001001001, 32'b00111110111100010000101110100101, 32'b00111110111100010100000100100100, 32'b00111110111100010111011011000110, 32'b00111110111100011010110010001101, 32'b00111110111100011110001001110111, 32'b00111110111100100001100010000110, 32'b00111110111100100100111010111001, 32'b00111110111100101000010100010000, 32'b00111110111100101011101110001100, 32'b00111110111100101111001000101101, 32'b00111110111100110010100011110011, 32'b00111110111100110101111111011110, 32'b00111110111100111001011011101110, 32'b00111110111100111100111000100011, 32'b00111110111101000000010101111111, 32'b00111110111101000011110100000000, 32'b00111110111101000111010010100111, 32'b00111110111101001010110001110100, 32'b00111110111101001110010001100111, 32'b00111110111101010001110010000001, 32'b00111110111101010101010011000001, 32'b00111110111101011000110100101000, 32'b00111110111101011100010110110110, 32'b00111110111101011111111001101100, 32'b00111110111101100011011101001000, 32'b00111110111101100111000001001100, 32'b00111110111101101010100101111000, 32'b00111110111101101110001011001100, 32'b00111110111101110001110001001000, 32'b00111110111101110101010111101100, 32'b00111110111101111000111110111000, 32'b00111110111101111100100110101101, 32'b00111110111110000000001111001011, 32'b00111110111110000011111000010001, 32'b00111110111110000111100010000001, 32'b00111110111110001011001100011010, 32'b00111110111110001110110111011101, 32'b00111110111110010010100011001001, 32'b00111110111110010110001111100000, 32'b00111110111110011001111100100000, 32'b00111110111110011101101010001011, 32'b00111110111110100001011000100000, 32'b00111110111110100101000111100000, 32'b00111110111110101000110111001011, 32'b00111110111110101100100111100001, 32'b00111110111110110000011000100011, 32'b00111110111110110100001010010000, 32'b00111110111110110111111100101000, 32'b00111110111110111011101111101101, 32'b00111110111110111111100011011101, 32'b00111110111111000011010111111010, 32'b00111110111111000111001101000100, 32'b00111110111111001011000010111010, 32'b00111110111111001110111001011101, 32'b00111110111111010010110000101110, 32'b00111110111111010110101000101011, 32'b00111110111111011010100001010111, 32'b00111110111111011110011010110000, 32'b00111110111111100010010100111000, 32'b00111110111111100110001111101101, 32'b00111110111111101010001011010010, 32'b00111110111111101110000111100100, 32'b00111110111111110010000100100110, 32'b00111110111111110110000010010111, 32'b00111110111111111010000000111000, 32'b00111110111111111110000000001000};
    assign b_table = '{32'b00111111100001011100001111001101, 32'b00111111100001011011000110100111, 32'b00111111100001011001111101111110, 32'b00111111100001011000110101010010, 32'b00111111100001010111101100100100, 32'b00111111100001010110100011110100, 32'b00111111100001010101011011000001, 32'b00111111100001010100010010001011, 32'b00111111100001010011001001010100, 32'b00111111100001010010000000011001, 32'b00111111100001010000110111011100, 32'b00111111100001001111101110011101, 32'b00111111100001001110100101011011, 32'b00111111100001001101011100010111, 32'b00111111100001001100010011010000, 32'b00111111100001001011001010000110, 32'b00111111100001001010000000111010, 32'b00111111100001001000110111101100, 32'b00111111100001000111101110011011, 32'b00111111100001000110100101000111, 32'b00111111100001000101011011110001, 32'b00111111100001000100010010011001, 32'b00111111100001000011001000111110, 32'b00111111100001000001111111100000, 32'b00111111100001000000110110000000, 32'b00111111100000111111101100011101, 32'b00111111100000111110100010110111, 32'b00111111100000111101011001010000, 32'b00111111100000111100001111100101, 32'b00111111100000111011000101111000, 32'b00111111100000111001111100001000, 32'b00111111100000111000110010010110, 32'b00111111100000110111101000100001, 32'b00111111100000110110011110101010, 32'b00111111100000110101010100110000, 32'b00111111100000110100001010110011, 32'b00111111100000110011000000110100, 32'b00111111100000110001110110110010, 32'b00111111100000110000101100101110, 32'b00111111100000101111100010100110, 32'b00111111100000101110011000011101, 32'b00111111100000101101001110010000, 32'b00111111100000101100000100000001, 32'b00111111100000101010111001110000, 32'b00111111100000101001101111011100, 32'b00111111100000101000100101000101, 32'b00111111100000100111011010101011, 32'b00111111100000100110010000001111, 32'b00111111100000100101000101110000, 32'b00111111100000100011111011001111, 32'b00111111100000100010110000101011, 32'b00111111100000100001100110000100, 32'b00111111100000100000011011011010, 32'b00111111100000011111010000101110, 32'b00111111100000011110000101111111, 32'b00111111100000011100111011001110, 32'b00111111100000011011110000011001, 32'b00111111100000011010100101100010, 32'b00111111100000011001011010101001, 32'b00111111100000011000001111101100, 32'b00111111100000010111000100101101, 32'b00111111100000010101111001101011, 32'b00111111100000010100101110100111, 32'b00111111100000010011100011100000, 32'b00111111100000010010011000010110, 32'b00111111100000010001001101001001, 32'b00111111100000010000000001111010, 32'b00111111100000001110110110100111, 32'b00111111100000001101101011010010, 32'b00111111100000001100011111111011, 32'b00111111100000001011010100100000, 32'b00111111100000001010001001000011, 32'b00111111100000001000111101100011, 32'b00111111100000000111110010000000, 32'b00111111100000000110100110011011, 32'b00111111100000000101011010110011, 32'b00111111100000000100001111000111, 32'b00111111100000000011000011011010, 32'b00111111100000000001110111101001, 32'b00111111100000000000101011110101, 32'b00111111011111111110111111111110, 32'b00111111011111111100101000001100, 32'b00111111011111111010010000010100, 32'b00111111011111110111111000010111, 32'b00111111011111110101100000010011, 32'b00111111011111110011001000001011, 32'b00111111011111110000101111111100, 32'b00111111011111101110010111101000, 32'b00111111011111101011111111001110, 32'b00111111011111101001100110101110, 32'b00111111011111100111001110001001, 32'b00111111011111100100110101011110, 32'b00111111011111100010011100101101, 32'b00111111011111100000000011110111, 32'b00111111011111011101101010111011, 32'b00111111011111011011010001111001, 32'b00111111011111011000111000110001, 32'b00111111011111010110011111100100, 32'b00111111011111010100000110010000, 32'b00111111011111010001101100110111, 32'b00111111011111001111010011011000, 32'b00111111011111001100111001110011, 32'b00111111011111001010100000001001, 32'b00111111011111001000000110011000, 32'b00111111011111000101101100100010, 32'b00111111011111000011010010100110, 32'b00111111011111000000111000100100, 32'b00111111011110111110011110011100, 32'b00111111011110111100000100001110, 32'b00111111011110111001101001111010, 32'b00111111011110110111001111100001, 32'b00111111011110110100110101000001, 32'b00111111011110110010011010011011, 32'b00111111011110101111111111110000, 32'b00111111011110101101100100111111, 32'b00111111011110101011001010000111, 32'b00111111011110101000101111001010, 32'b00111111011110100110010100000110, 32'b00111111011110100011111000111101, 32'b00111111011110100001011101101110, 32'b00111111011110011111000010011000, 32'b00111111011110011100100110111101, 32'b00111111011110011010001011011011, 32'b00111111011110010111101111110100, 32'b00111111011110010101010100000110, 32'b00111111011110010010111000010010, 32'b00111111011110010000011100011000, 32'b00111111011110001110000000011000, 32'b00111111011110001011100100010010, 32'b00111111011110001001001000000110, 32'b00111111011110000110101011110100, 32'b00111111011110000100001111011011, 32'b00111111011110000001110010111101, 32'b00111111011101111111010110011000, 32'b00111111011101111100111001101101, 32'b00111111011101111010011100111100, 32'b00111111011101111000000000000101, 32'b00111111011101110101100011000111, 32'b00111111011101110011000110000011, 32'b00111111011101110000101000111001, 32'b00111111011101101110001011101001, 32'b00111111011101101011101110010010, 32'b00111111011101101001010000110101, 32'b00111111011101100110110011010010, 32'b00111111011101100100010101101001, 32'b00111111011101100001110111111001, 32'b00111111011101011111011010000011, 32'b00111111011101011100111100000111, 32'b00111111011101011010011110000100, 32'b00111111011101010111111111111011, 32'b00111111011101010101100001101011, 32'b00111111011101010011000011010101, 32'b00111111011101010000100100111001, 32'b00111111011101001110000110010110, 32'b00111111011101001011100111101101, 32'b00111111011101001001001000111110, 32'b00111111011101000110101010001000, 32'b00111111011101000100001011001011, 32'b00111111011101000001101100001001, 32'b00111111011100111111001100111111, 32'b00111111011100111100101101101111, 32'b00111111011100111010001110011001, 32'b00111111011100110111101110111100, 32'b00111111011100110101001111011001, 32'b00111111011100110010101111101111, 32'b00111111011100110000001111111110, 32'b00111111011100101101110000000111, 32'b00111111011100101011010000001001, 32'b00111111011100101000110000000101, 32'b00111111011100100110001111111010, 32'b00111111011100100011101111101001, 32'b00111111011100100001001111010001, 32'b00111111011100011110101110110010, 32'b00111111011100011100001110001101, 32'b00111111011100011001101101100000, 32'b00111111011100010111001100101110, 32'b00111111011100010100101011110100, 32'b00111111011100010010001010110100, 32'b00111111011100001111101001101101, 32'b00111111011100001101001000011111, 32'b00111111011100001010100111001011, 32'b00111111011100001000000101110000, 32'b00111111011100000101100100001110, 32'b00111111011100000011000010100101, 32'b00111111011100000000100000110110, 32'b00111111011011111101111110111111, 32'b00111111011011111011011101000010, 32'b00111111011011111000111010111110, 32'b00111111011011110110011000110011, 32'b00111111011011110011110110100010, 32'b00111111011011110001010100001001, 32'b00111111011011101110110001101010, 32'b00111111011011101100001111000011, 32'b00111111011011101001101100010110, 32'b00111111011011100111001001100001, 32'b00111111011011100100100110100110, 32'b00111111011011100010000011100100, 32'b00111111011011011111100000011011, 32'b00111111011011011100111101001011, 32'b00111111011011011010011001110011, 32'b00111111011011010111110110010101, 32'b00111111011011010101010010110000, 32'b00111111011011010010101111000100, 32'b00111111011011010000001011010000, 32'b00111111011011001101100111010110, 32'b00111111011011001011000011010100, 32'b00111111011011001000011111001100, 32'b00111111011011000101111010111100, 32'b00111111011011000011010110100101, 32'b00111111011011000000110010000111, 32'b00111111011010111110001101100010, 32'b00111111011010111011101000110101, 32'b00111111011010111001000100000010, 32'b00111111011010110110011111000111, 32'b00111111011010110011111010000101, 32'b00111111011010110001010100111011, 32'b00111111011010101110101111101011, 32'b00111111011010101100001010010011, 32'b00111111011010101001100100110100, 32'b00111111011010100110111111001101, 32'b00111111011010100100011001100000, 32'b00111111011010100001110011101011, 32'b00111111011010011111001101101110, 32'b00111111011010011100100111101010, 32'b00111111011010011010000001011111, 32'b00111111011010010111011011001101, 32'b00111111011010010100110100110011, 32'b00111111011010010010001110010001, 32'b00111111011010001111100111101001, 32'b00111111011010001101000000111000, 32'b00111111011010001010011010000001, 32'b00111111011010000111110011000001, 32'b00111111011010000101001011111011, 32'b00111111011010000010100100101100, 32'b00111111011001111111111101010111, 32'b00111111011001111101010101111001, 32'b00111111011001111010101110010101, 32'b00111111011001111000000110101000, 32'b00111111011001110101011110110100, 32'b00111111011001110010110110111000, 32'b00111111011001110000001110110101, 32'b00111111011001101101100110101010, 32'b00111111011001101010111110010111, 32'b00111111011001101000010101111101, 32'b00111111011001100101101101011011, 32'b00111111011001100011000100110001, 32'b00111111011001100000011100000000, 32'b00111111011001011101110011000111, 32'b00111111011001011011001010000110, 32'b00111111011001011000100000111101, 32'b00111111011001010101110111101101, 32'b00111111011001010011001110010100, 32'b00111111011001010000100100110100, 32'b00111111011001001101111011001100, 32'b00111111011001001011010001011100, 32'b00111111011001001000100111100101, 32'b00111111011001000101111101100101, 32'b00111111011001000011010011011101, 32'b00111111011001000000101001001110, 32'b00111111011000111101111110110111, 32'b00111111011000111011010100010111, 32'b00111111011000111000101001110000, 32'b00111111011000110101111111000000, 32'b00111111011000110011010100001001, 32'b00111111011000110000101001001010, 32'b00111111011000101101111110000010, 32'b00111111011000101011010010110010, 32'b00111111011000101000100111011011, 32'b00111111011000100101111011111011, 32'b00111111011000100011010000010011, 32'b00111111011000100000100100100011, 32'b00111111011000011101111000101011, 32'b00111111011000011011001100101011, 32'b00111111011000011000100000100010, 32'b00111111011000010101110100010001, 32'b00111111011000010011000111111000, 32'b00111111011000010000011011010111, 32'b00111111011000001101101110101101, 32'b00111111011000001011000001111011, 32'b00111111011000001000010101000001, 32'b00111111011000000101100111111111, 32'b00111111011000000010111010110100, 32'b00111111011000000000001101100001, 32'b00111111010111111101100000000101, 32'b00111111010111111010110010100001, 32'b00111111010111111000000100110101, 32'b00111111010111110101010111000000, 32'b00111111010111110010101001000011, 32'b00111111010111101111111010111101, 32'b00111111010111101101001100101110, 32'b00111111010111101010011110011000, 32'b00111111010111100111101111111000, 32'b00111111010111100101000001010000, 32'b00111111010111100010010010100000, 32'b00111111010111011111100011100111, 32'b00111111010111011100110100100101, 32'b00111111010111011010000101011011, 32'b00111111010111010111010110001000, 32'b00111111010111010100100110101100, 32'b00111111010111010001110111001000, 32'b00111111010111001111000111011010, 32'b00111111010111001100010111100101, 32'b00111111010111001001100111100110, 32'b00111111010111000110110111011111, 32'b00111111010111000100000111001110, 32'b00111111010111000001010110110101, 32'b00111111010110111110100110010011, 32'b00111111010110111011110101101001, 32'b00111111010110111001000100110101, 32'b00111111010110110110010011111001, 32'b00111111010110110011100010110011, 32'b00111111010110110000110001100101, 32'b00111111010110101110000000001101, 32'b00111111010110101011001110101101, 32'b00111111010110101000011101000100, 32'b00111111010110100101101011010001, 32'b00111111010110100010111001010110, 32'b00111111010110100000000111010001, 32'b00111111010110011101010101000100, 32'b00111111010110011010100010101101, 32'b00111111010110010111110000001101, 32'b00111111010110010100111101100100, 32'b00111111010110010010001010110010, 32'b00111111010110001111010111110110, 32'b00111111010110001100100100110010, 32'b00111111010110001001110001100100, 32'b00111111010110000110111110001101, 32'b00111111010110000100001010101100, 32'b00111111010110000001010111000010, 32'b00111111010101111110100011001111, 32'b00111111010101111011101111010011, 32'b00111111010101111000111011001101, 32'b00111111010101110110000110111101, 32'b00111111010101110011010010100101, 32'b00111111010101110000011110000010, 32'b00111111010101101101101001010111, 32'b00111111010101101010110100100001, 32'b00111111010101100111111111100011, 32'b00111111010101100101001010011010, 32'b00111111010101100010010101001001, 32'b00111111010101011111011111101101, 32'b00111111010101011100101010001000, 32'b00111111010101011001110100011001, 32'b00111111010101010110111110100001, 32'b00111111010101010100001000011111, 32'b00111111010101010001010010010011, 32'b00111111010101001110011011111101, 32'b00111111010101001011100101011110, 32'b00111111010101001000101110110101, 32'b00111111010101000101111000000010, 32'b00111111010101000011000001000101, 32'b00111111010101000000001001111111, 32'b00111111010100111101010010101110, 32'b00111111010100111010011011010100, 32'b00111111010100110111100011101111, 32'b00111111010100110100101100000001, 32'b00111111010100110001110100001001, 32'b00111111010100101110111100000110, 32'b00111111010100101100000011111010, 32'b00111111010100101001001011100011, 32'b00111111010100100110010011000011, 32'b00111111010100100011011010011000, 32'b00111111010100100000100001100011, 32'b00111111010100011101101000100100, 32'b00111111010100011010101111011011, 32'b00111111010100010111110110000111, 32'b00111111010100010100111100101010, 32'b00111111010100010010000011000010, 32'b00111111010100001111001001001111, 32'b00111111010100001100001111010011, 32'b00111111010100001001010101001100, 32'b00111111010100000110011010111010, 32'b00111111010100000011100000011111, 32'b00111111010100000000100101111000, 32'b00111111010011111101101011001000, 32'b00111111010011111010110000001101, 32'b00111111010011110111110101000111, 32'b00111111010011110100111001110111, 32'b00111111010011110001111110011100, 32'b00111111010011101111000010110110, 32'b00111111010011101100000111000110, 32'b00111111010011101001001011001011, 32'b00111111010011100110001111000110, 32'b00111111010011100011010010110110, 32'b00111111010011100000010110011011, 32'b00111111010011011101011001110101, 32'b00111111010011011010011101000100, 32'b00111111010011010111100000001001, 32'b00111111010011010100100011000011, 32'b00111111010011010001100101110010, 32'b00111111010011001110101000010110, 32'b00111111010011001011101010101111, 32'b00111111010011001000101100111101, 32'b00111111010011000101101111000000, 32'b00111111010011000010110000111000, 32'b00111111010010111111110010100101, 32'b00111111010010111100110100000110, 32'b00111111010010111001110101011101, 32'b00111111010010110110110110101000, 32'b00111111010010110011110111101001, 32'b00111111010010110000111000011110, 32'b00111111010010101101111001000111, 32'b00111111010010101010111001100110, 32'b00111111010010100111111001111001, 32'b00111111010010100100111010000001, 32'b00111111010010100001111001111101, 32'b00111111010010011110111001101110, 32'b00111111010010011011111001010100, 32'b00111111010010011000111000101110, 32'b00111111010010010101110111111101, 32'b00111111010010010010110111000000, 32'b00111111010010001111110101110111, 32'b00111111010010001100110100100011, 32'b00111111010010001001110011000011, 32'b00111111010010000110110001011000, 32'b00111111010010000011101111100000, 32'b00111111010010000000101101011101, 32'b00111111010001111101101011001111, 32'b00111111010001111010101000110100, 32'b00111111010001110111100110001110, 32'b00111111010001110100100011011100, 32'b00111111010001110001100000011101, 32'b00111111010001101110011101010011, 32'b00111111010001101011011001111101, 32'b00111111010001101000010110011011, 32'b00111111010001100101010010101101, 32'b00111111010001100010001110110011, 32'b00111111010001011111001010101101, 32'b00111111010001011100000110011010, 32'b00111111010001011001000001111011, 32'b00111111010001010101111101010000, 32'b00111111010001010010111000011001, 32'b00111111010001001111110011010110, 32'b00111111010001001100101110000110, 32'b00111111010001001001101000101010, 32'b00111111010001000110100011000001, 32'b00111111010001000011011101001100, 32'b00111111010001000000010111001011, 32'b00111111010000111101010000111101, 32'b00111111010000111010001010100010, 32'b00111111010000110111000011111011, 32'b00111111010000110011111101000111, 32'b00111111010000110000110110000111, 32'b00111111010000101101101110111010, 32'b00111111010000101010100111100000, 32'b00111111010000100111011111111001, 32'b00111111010000100100011000000110, 32'b00111111010000100001010000000110, 32'b00111111010000011110000111111000, 32'b00111111010000011010111111011110, 32'b00111111010000010111110110110111, 32'b00111111010000010100101110000011, 32'b00111111010000010001100101000010, 32'b00111111010000001110011011110011, 32'b00111111010000001011010010011000, 32'b00111111010000001000001000101111, 32'b00111111010000000100111110111010, 32'b00111111010000000001110100110111, 32'b00111111001111111110101010100110, 32'b00111111001111111011100000001000, 32'b00111111001111111000010101011101, 32'b00111111001111110101001010100101, 32'b00111111001111110001111111011111, 32'b00111111001111101110110100001100, 32'b00111111001111101011101000101011, 32'b00111111001111101000011100111100, 32'b00111111001111100101010001000000, 32'b00111111001111100010000100110110, 32'b00111111001111011110111000011110, 32'b00111111001111011011101011111001, 32'b00111111001111011000011111000110, 32'b00111111001111010101010010000101, 32'b00111111001111010010000100110110, 32'b00111111001111001110110111011001, 32'b00111111001111001011101001101110, 32'b00111111001111001000011011110101, 32'b00111111001111000101001101101110, 32'b00111111001111000001111111011001, 32'b00111111001110111110110000110110, 32'b00111111001110111011100010000101, 32'b00111111001110111000010011000101, 32'b00111111001110110101000011110111, 32'b00111111001110110001110100011011, 32'b00111111001110101110100100110000, 32'b00111111001110101011010100110111, 32'b00111111001110101000000100110000, 32'b00111111001110100100110100011010, 32'b00111111001110100001100011110101, 32'b00111111001110011110010011000010, 32'b00111111001110011011000010000000, 32'b00111111001110010111110000101111, 32'b00111111001110010100011111010000, 32'b00111111001110010001001101100001, 32'b00111111001110001101111011100100, 32'b00111111001110001010101001011000, 32'b00111111001110000111010110111101, 32'b00111111001110000100000100010011, 32'b00111111001110000000110001011010, 32'b00111111001101111101011110010010, 32'b00111111001101111010001010111010, 32'b00111111001101110110110111010011, 32'b00111111001101110011100011011110, 32'b00111111001101110000001111011000, 32'b00111111001101101100111011000100, 32'b00111111001101101001100110100000, 32'b00111111001101100110010001101100, 32'b00111111001101100010111100101001, 32'b00111111001101011111100111010110, 32'b00111111001101011100010001110100, 32'b00111111001101011000111100000010, 32'b00111111001101010101100110000000, 32'b00111111001101010010001111101111, 32'b00111111001101001111100110100010, 32'b00111111001101001110001011111110, 32'b00111111001101001100110001011000, 32'b00111111001101001011010110101111, 32'b00111111001101001001111100000011, 32'b00111111001101001000100001010100, 32'b00111111001101000111000110100011, 32'b00111111001101000101101011101110, 32'b00111111001101000100010000110111, 32'b00111111001101000010110101111100, 32'b00111111001101000001011010111111, 32'b00111111001100111111111111111111, 32'b00111111001100111110100100111100, 32'b00111111001100111101001001110111, 32'b00111111001100111011101110101110, 32'b00111111001100111010010011100011, 32'b00111111001100111000111000010100, 32'b00111111001100110111011101000011, 32'b00111111001100110110000001101111, 32'b00111111001100110100100110010111, 32'b00111111001100110011001010111101, 32'b00111111001100110001101111100000, 32'b00111111001100110000010100000001, 32'b00111111001100101110111000011110, 32'b00111111001100101101011100111000, 32'b00111111001100101100000001001111, 32'b00111111001100101010100101100100, 32'b00111111001100101001001001110101, 32'b00111111001100100111101110000100, 32'b00111111001100100110010010001111, 32'b00111111001100100100110110011000, 32'b00111111001100100011011010011110, 32'b00111111001100100001111110100000, 32'b00111111001100100000100010100000, 32'b00111111001100011111000110011101, 32'b00111111001100011101101010010111, 32'b00111111001100011100001110001101, 32'b00111111001100011010110010000001, 32'b00111111001100011001010101110010, 32'b00111111001100010111111001100000, 32'b00111111001100010110011101001011, 32'b00111111001100010101000000110011, 32'b00111111001100010011100100010111, 32'b00111111001100010010000111111001, 32'b00111111001100010000101011011000, 32'b00111111001100001111001110110100, 32'b00111111001100001101110010001100, 32'b00111111001100001100010101100010, 32'b00111111001100001010111000110101, 32'b00111111001100001001011100000100, 32'b00111111001100000111111111010001, 32'b00111111001100000110100010011010, 32'b00111111001100000101000101100001, 32'b00111111001100000011101000100100, 32'b00111111001100000010001011100101, 32'b00111111001100000000101110100010, 32'b00111111001011111111010001011100, 32'b00111111001011111101110100010011, 32'b00111111001011111100010111000111, 32'b00111111001011111010111001111000, 32'b00111111001011111001011100100110, 32'b00111111001011110111111111010001, 32'b00111111001011110110100001111000, 32'b00111111001011110101000100011101, 32'b00111111001011110011100110111110, 32'b00111111001011110010001001011100, 32'b00111111001011110000101011111000, 32'b00111111001011101111001110010000, 32'b00111111001011101101110000100101, 32'b00111111001011101100010010110110, 32'b00111111001011101010110101000101, 32'b00111111001011101001010111010000, 32'b00111111001011100111111001011001, 32'b00111111001011100110011011011110, 32'b00111111001011100100111101100000, 32'b00111111001011100011011111011111, 32'b00111111001011100010000001011010, 32'b00111111001011100000100011010011, 32'b00111111001011011111000101001000, 32'b00111111001011011101100110111010, 32'b00111111001011011100001000101001, 32'b00111111001011011010101010010101, 32'b00111111001011011001001011111101, 32'b00111111001011010111101101100011, 32'b00111111001011010110001111000101, 32'b00111111001011010100110000100100, 32'b00111111001011010011010001111111, 32'b00111111001011010001110011011000, 32'b00111111001011010000010100101101, 32'b00111111001011001110110101111111, 32'b00111111001011001101010111001110, 32'b00111111001011001011111000011001, 32'b00111111001011001010011001100001, 32'b00111111001011001000111010100110, 32'b00111111001011000111011011101000, 32'b00111111001011000101111100100110, 32'b00111111001011000100011101100001, 32'b00111111001011000010111110011001, 32'b00111111001011000001011111001110, 32'b00111111001010111111111111111111, 32'b00111111001010111110100000101101, 32'b00111111001010111101000001011000, 32'b00111111001010111011100001111111, 32'b00111111001010111010000010100011, 32'b00111111001010111000100011000100, 32'b00111111001010110111000011100001, 32'b00111111001010110101100011111011, 32'b00111111001010110100000100010010, 32'b00111111001010110010100100100110, 32'b00111111001010110001000100110110, 32'b00111111001010101111100101000010, 32'b00111111001010101110000101001100, 32'b00111111001010101100100101010010, 32'b00111111001010101011000101010100, 32'b00111111001010101001100101010100, 32'b00111111001010101000000101001111, 32'b00111111001010100110100101001000, 32'b00111111001010100101000100111101, 32'b00111111001010100011100100101111, 32'b00111111001010100010000100011101, 32'b00111111001010100000100100001000, 32'b00111111001010011111000011101111, 32'b00111111001010011101100011010011, 32'b00111111001010011100000010110100, 32'b00111111001010011010100010010001, 32'b00111111001010011001000001101011, 32'b00111111001010010111100001000001, 32'b00111111001010010110000000010100, 32'b00111111001010010100011111100100, 32'b00111111001010010010111110110000, 32'b00111111001010010001011101111000, 32'b00111111001010001111111100111101, 32'b00111111001010001110011011111111, 32'b00111111001010001100111010111101, 32'b00111111001010001011011001110111, 32'b00111111001010001001111000101111, 32'b00111111001010001000010111100010, 32'b00111111001010000110110110010010, 32'b00111111001010000101010100111111, 32'b00111111001010000011110011101000, 32'b00111111001010000010010010001101, 32'b00111111001010000000110000101111, 32'b00111111001001111111001111001110, 32'b00111111001001111101101101101001, 32'b00111111001001111100001100000000, 32'b00111111001001111010101010010100, 32'b00111111001001111001001000100100, 32'b00111111001001110111100110110001, 32'b00111111001001110110000100111010, 32'b00111111001001110100100011000000, 32'b00111111001001110011000001000010, 32'b00111111001001110001011111000000, 32'b00111111001001101111111100111011, 32'b00111111001001101110011010110010, 32'b00111111001001101100111000100110, 32'b00111111001001101011010110010110, 32'b00111111001001101001110100000010, 32'b00111111001001101000010001101011, 32'b00111111001001100110101111010000, 32'b00111111001001100101001100110001, 32'b00111111001001100011101010001111, 32'b00111111001001100010000111101001, 32'b00111111001001100000100101000000, 32'b00111111001001011111000010010010, 32'b00111111001001011101011111100010, 32'b00111111001001011011111100101101, 32'b00111111001001011010011001110101, 32'b00111111001001011000110110111001, 32'b00111111001001010111010011111001, 32'b00111111001001010101110000110110, 32'b00111111001001010100001101101111, 32'b00111111001001010010101010100100, 32'b00111111001001010001000111010110, 32'b00111111001001001111100100000100, 32'b00111111001001001110000000101110, 32'b00111111001001001100011101010100, 32'b00111111001001001010111001110111, 32'b00111111001001001001010110010101, 32'b00111111001001000111110010110000, 32'b00111111001001000110001111001000, 32'b00111111001001000100101011011011, 32'b00111111001001000011000111101011, 32'b00111111001001000001100011110111, 32'b00111111001000111111111111111111, 32'b00111111001000111110011100000011, 32'b00111111001000111100111000000100, 32'b00111111001000111011010100000001, 32'b00111111001000111001101111111010, 32'b00111111001000111000001011101111, 32'b00111111001000110110100111100000, 32'b00111111001000110101000011001101, 32'b00111111001000110011011110110111, 32'b00111111001000110001111010011100, 32'b00111111001000110000010101111110, 32'b00111111001000101110110001011100, 32'b00111111001000101101001100110110, 32'b00111111001000101011101000001100, 32'b00111111001000101010000011011111, 32'b00111111001000101000011110101101, 32'b00111111001000100110111001110111, 32'b00111111001000100101010100111110, 32'b00111111001000100011110000000001, 32'b00111111001000100010001010111111, 32'b00111111001000100000100101111010, 32'b00111111001000011111000000110001, 32'b00111111001000011101011011100100, 32'b00111111001000011011110110010011, 32'b00111111001000011010010000111110, 32'b00111111001000011000101011100100, 32'b00111111001000010111000110000111, 32'b00111111001000010101100000100110, 32'b00111111001000010011111011000001, 32'b00111111001000010010010101011000, 32'b00111111001000010000101111101011, 32'b00111111001000001111001001111010, 32'b00111111001000001101100100000101, 32'b00111111001000001011111110001100, 32'b00111111001000001010011000001111, 32'b00111111001000001000110010001110, 32'b00111111001000000111001100001001, 32'b00111111001000000101100110000000, 32'b00111111001000000011111111110010, 32'b00111111001000000010011001100001, 32'b00111111001000000000110011001011, 32'b00111111000111111111001100110010, 32'b00111111000111111101100110010100, 32'b00111111000111111011111111110010, 32'b00111111000111111010011001001100, 32'b00111111000111111000110010100010, 32'b00111111000111110111001011110100, 32'b00111111000111110101100101000010, 32'b00111111000111110011111110001011, 32'b00111111000111110010010111010001, 32'b00111111000111110000110000010010, 32'b00111111000111101111001001001111, 32'b00111111000111101101100010001000, 32'b00111111000111101011111010111100, 32'b00111111000111101010010011101101, 32'b00111111000111101000101100011001, 32'b00111111000111100111000101000001, 32'b00111111000111100101011101100101, 32'b00111111000111100011110110000101, 32'b00111111000111100010001110100000, 32'b00111111000111100000100110110111, 32'b00111111000111011110111111001010, 32'b00111111000111011101010111011001, 32'b00111111000111011011101111100011, 32'b00111111000111011010000111101001, 32'b00111111000111011000011111101011, 32'b00111111000111010110110111101001, 32'b00111111000111010101001111100010, 32'b00111111000111010011100111010111, 32'b00111111000111010001111111001000, 32'b00111111000111010000010110110100, 32'b00111111000111001110101110011100, 32'b00111111000111001101000101111111, 32'b00111111000111001011011101011111, 32'b00111111000111001001110100111010, 32'b00111111000111001000001100010000, 32'b00111111000111000110100011100010, 32'b00111111000111000100111010110000, 32'b00111111000111000011010001111001, 32'b00111111000111000001101000111110, 32'b00111111000110111111111111111111, 32'b00111111000110111110010110111011, 32'b00111111000110111100101101110011, 32'b00111111000110111011000100100110, 32'b00111111000110111001011011010101, 32'b00111111000110110111110001111111, 32'b00111111000110110110001000100101, 32'b00111111000110110100011111000111, 32'b00111111000110110010110101100100, 32'b00111111000110110001001011111100, 32'b00111111000110101111100010010000, 32'b00111111000110101101111000100000, 32'b00111111000110101100001110101010, 32'b00111111000110101010100100110001, 32'b00111111000110101000111010110011, 32'b00111111000110100111010000110000, 32'b00111111000110100101100110101001, 32'b00111111000110100011111100011101, 32'b00111111000110100010010010001101, 32'b00111111000110100000100111111000, 32'b00111111000110011110111101011110, 32'b00111111000110011101010011000000, 32'b00111111000110011011101000011110, 32'b00111111000110011001111101110110, 32'b00111111000110011000010011001010, 32'b00111111000110010110101000011010, 32'b00111111000110010100111101100100, 32'b00111111000110010011010010101010, 32'b00111111000110010001100111101100, 32'b00111111000110001111111100101001, 32'b00111111000110001110010001100001, 32'b00111111000110001100100110010100, 32'b00111111000110001010111011000011, 32'b00111111000110001001001111101101, 32'b00111111000110000111100100010010, 32'b00111111000110000101111000110010, 32'b00111111000110000100001101001110, 32'b00111111000110000010100001100101, 32'b00111111000110000000110101110111, 32'b00111111000101111111001010000101, 32'b00111111000101111101011110001110, 32'b00111111000101111011110010010010, 32'b00111111000101111010000110010001, 32'b00111111000101111000011010001011, 32'b00111111000101110110101110000000, 32'b00111111000101110101000001110001, 32'b00111111000101110011010101011101, 32'b00111111000101110001101001000100, 32'b00111111000101101111111100100110, 32'b00111111000101101110010000000011, 32'b00111111000101101100100011011011, 32'b00111111000101101010110110101111, 32'b00111111000101101001001001111101, 32'b00111111000101100111011101000111, 32'b00111111000101100101110000001011, 32'b00111111000101100100000011001011, 32'b00111111000101100010010110000110, 32'b00111111000101100000101000111100, 32'b00111111000101011110111011101101, 32'b00111111000101011101001110011001, 32'b00111111000101011011100001000000, 32'b00111111000101011001110011100001, 32'b00111111000101011000000101111110, 32'b00111111000101010110011000010110, 32'b00111111000101010100101010101001, 32'b00111111000101010010111100110111, 32'b00111111000101010001001111000000, 32'b00111111000101001111100001000011, 32'b00111111000101001101110011000010, 32'b00111111000101001100000100111011, 32'b00111111000101001010010110110000, 32'b00111111000101001000101000011111, 32'b00111111000101000110111010001001, 32'b00111111000101000101001011101110, 32'b00111111000101000011011101001110, 32'b00111111000101000001101110101001, 32'b00111111000100111111111111111111, 32'b00111111000100111110010001001111, 32'b00111111000100111100100010011010, 32'b00111111000100111010110011100000, 32'b00111111000100111001000100100001, 32'b00111111000100110111010101011101, 32'b00111111000100110101100110010011, 32'b00111111000100110011110111000100, 32'b00111111000100110010000111110000, 32'b00111111000100110000011000010111, 32'b00111111000100101110101000111000, 32'b00111111000100101100111001010100, 32'b00111111000100101011001001101011, 32'b00111111000100101001011001111101, 32'b00111111000100100111101010001001, 32'b00111111000100100101111010001111, 32'b00111111000100100100001010010001, 32'b00111111000100100010011010001101, 32'b00111111000100100000101010000100, 32'b00111111000100011110111001110101, 32'b00111111000100011101001001100001, 32'b00111111000100011011011001000111, 32'b00111111000100011001101000101000, 32'b00111111000100010111111000000100, 32'b00111111000100010110000111011010, 32'b00111111000100010100010110101011, 32'b00111111000100010010100101110110, 32'b00111111000100010000110100111100, 32'b00111111000100001111000011111100, 32'b00111111000100001101010010110111, 32'b00111111000100001011100001101100, 32'b00111111000100001001110000011100, 32'b00111111000100000111111111000110, 32'b00111111000100000110001101101011, 32'b00111111000100000100011100001010, 32'b00111111000100000010101010100011, 32'b00111111000100000000111000110111, 32'b00111111000011111111000111000101, 32'b00111111000011111101010101001110, 32'b00111111000011111011100011010001, 32'b00111111000011111001110001001110, 32'b00111111000011110111111111000101, 32'b00111111000011110110001100110111, 32'b00111111000011110100011010100100, 32'b00111111000011110010101000001010, 32'b00111111000011110000110101101011, 32'b00111111000011101111000011000110, 32'b00111111000011101101010000011100, 32'b00111111000011101011011101101011, 32'b00111111000011101001101010110101, 32'b00111111000011100111110111111001, 32'b00111111000011100110000100110111, 32'b00111111000011100100010001110000, 32'b00111111000011100010011110100010, 32'b00111111000011100000101011001111, 32'b00111111000011011110110111110110, 32'b00111111000011011101000100010111, 32'b00111111000011011011010000110010, 32'b00111111000011011001011101001000, 32'b00111111000011010111101001010111, 32'b00111111000011010101110101100000, 32'b00111111000011010100000001100100, 32'b00111111000011010010001101100010, 32'b00111111000011010000011001011001, 32'b00111111000011001110100101001011, 32'b00111111000011001100110000110110, 32'b00111111000011001010111100011100, 32'b00111111000011001001000111111100, 32'b00111111000011000111010011010101, 32'b00111111000011000101011110101001, 32'b00111111000011000011101001110110, 32'b00111111000011000001110100111101, 32'b00111111000010111111111111111110, 32'b00111111000010111110001010111010, 32'b00111111000010111100010101101111, 32'b00111111000010111010100000011101, 32'b00111111000010111000101011000110, 32'b00111111000010110110110101101001, 32'b00111111000010110101000000000101, 32'b00111111000010110011001010011011, 32'b00111111000010110001010100101011, 32'b00111111000010101111011110110101, 32'b00111111000010101101101000111000, 32'b00111111000010101011110010110101, 32'b00111111000010101001111100101100, 32'b00111111000010101000000110011100, 32'b00111111000010100110010000000111, 32'b00111111000010100100011001101011, 32'b00111111000010100010100011001000, 32'b00111111000010100000101100011111, 32'b00111111000010011110110101110000, 32'b00111111000010011100111110111011, 32'b00111111000010011011000111111111, 32'b00111111000010011001010000111100, 32'b00111111000010010111011001110011, 32'b00111111000010010101100010100100, 32'b00111111000010010011101011001110, 32'b00111111000010010001110011110010, 32'b00111111000010001111111100001111, 32'b00111111000010001110000100100110, 32'b00111111000010001100001100110110, 32'b00111111000010001010010101000000, 32'b00111111000010001000011101000011, 32'b00111111000010000110100100111111, 32'b00111111000010000100101100110101, 32'b00111111000010000010110100100100, 32'b00111111000010000000111100001101, 32'b00111111000001111111000011101110, 32'b00111111000001111101001011001010, 32'b00111111000001111011010010011110, 32'b00111111000001111001011001101100, 32'b00111111000001110111100000110011, 32'b00111111000001110101100111110011, 32'b00111111000001110011101110101101, 32'b00111111000001110001110101100000, 32'b00111111000001101111111100001100, 32'b00111111000001101110000010110001, 32'b00111111000001101100001001001111, 32'b00111111000001101010001111100110, 32'b00111111000001101000010101110111, 32'b00111111000001100110011100000001, 32'b00111111000001100100100010000011, 32'b00111111000001100010100111111111, 32'b00111111000001100000101101110100, 32'b00111111000001011110110011100010, 32'b00111111000001011100111001001001, 32'b00111111000001011010111110101001, 32'b00111111000001011001000100000010, 32'b00111111000001010111001001010100, 32'b00111111000001010101001110011111, 32'b00111111000001010011010011100010, 32'b00111111000001010001011000011111, 32'b00111111000001001111011101010101, 32'b00111111000001001101100010000011, 32'b00111111000001001011100110101010, 32'b00111111000001001001101011001010, 32'b00111111000001000111101111100011, 32'b00111111000001000101110011110101, 32'b00111111000001000011110111111111, 32'b00111111000001000001111100000010, 32'b00111111000000111111111111111110, 32'b00111111000000111110000011110011, 32'b00111111000000111100000111100000, 32'b00111111000000111010001011000110, 32'b00111111000000111000001110100101, 32'b00111111000000110110010001111100, 32'b00111111000000110100010101001100, 32'b00111111000000110010011000010100, 32'b00111111000000110000011011010101, 32'b00111111000000101110011110001110, 32'b00111111000000101100100001000000, 32'b00111111000000101010100011101011, 32'b00111111000000101000100110001110, 32'b00111111000000100110101000101001, 32'b00111111000000100100101010111101, 32'b00111111000000100010101101001010, 32'b00111111000000100000101111001110, 32'b00111111000000011110110001001011, 32'b00111111000000011100110011000001, 32'b00111111000000011010110100101111, 32'b00111111000000011000110110010101, 32'b00111111000000010110110111110011, 32'b00111111000000010100111001001010, 32'b00111111000000010010111010011000, 32'b00111111000000010000111011011111, 32'b00111111000000001110111100011111, 32'b00111111000000001100111101010110, 32'b00111111000000001010111110000110, 32'b00111111000000001000111110101101, 32'b00111111000000000110111111001101, 32'b00111111000000000100111111100101, 32'b00111111000000000010111111110101, 32'b00111111000000000000111111111101};

    wire [9:0] key0;
    assign key0 = (x[23]==1)? {1'b0, x[22:14]} : {1'b1, x[22:14]};
    wire [7:0] y_sub_e0;
    assign y_sub_e0 = ((x[30:23]-8'd127)>>1)+8'd127;
    reg [9:0] key_1;
    reg [7:0] y_sub_e_1;
    reg [7:0] y_sub_e_2;
    reg [7:0] y_sub_e_3;
    reg [7:0] y_sub_e_4;
    reg [7:0] y_sub_e_5;
    reg [31:0] x1;
    reg [31:0] x2;
    reg [31:0] x3;
    reg [31:0] x4;
    reg [31:0] x5;
    always @(posedge clk) begin
        key_1 <= key0;
        y_sub_e_1 <= y_sub_e0;
        x1 <= x;
        x2 <= x1;
        x3 <= x2;
        x4 <= x3;
        x5 <= x4;
        
    end

    wire [31:0] ax3; 
    wire [31:0] test_a1;
    wire [31:0] test_b1;

    assign test_a1 = a_table[key_1];
    assign test_b1 = b_table[key_1];
    wire [31:0] x_m1;
    assign x_m1 = (x1[23]==1)?{1'b0, 8'd127, x1[22:0]}:{1'b0, 8'd128, x1[22:0]};
    fmul fmull(test_a1,x_m1,ax3,clk);
    reg [31:0] test_b_2;
    reg [31:0] test_b_3;


    always @(posedge clk) begin
        test_b_2 <= test_b1;
        test_b_3 <= test_b_2;
        y_sub_e_2 <= y_sub_e_1;
        y_sub_e_3 <= y_sub_e_2;
        y_sub_e_4 <= y_sub_e_3;
        y_sub_e_5 <= y_sub_e_4;
    end
    wire [31:0] y_sub5;
    fadd faddd(test_b_3,ax3,y_sub5,clk);
    wire [31:0] y_sub55;
    assign y_sub55 = {1'b0,y_sub_e_5, y_sub5[22:0] };
    assign y = (x5[31]==1) ? 32'b01111111100000000000000000000000 : y_sub55;

    

endmodule