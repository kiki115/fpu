`default_nettype none
`include "fadd.sv"
/* verilator lint_off MULTITOP */
// hi
module finv (input wire [31:0]  x,
             output wire [31:0] y,
            input wire clk);

    wire [31:0] a_table[1023:0];
    wire [31:0] b_table[1023:0];
    assign a_table = '{32'b10111110100000000001000000000010, 32'b10111110100000000011000000001110, 32'b10111110100000000101000000100110, 32'b10111110100000000111000001001010, 32'b10111110100000001001000001111010, 32'b10111110100000001011000010110111, 32'b10111110100000001101000011111111, 32'b10111110100000001111000101010100, 32'b10111110100000010001000110110100, 32'b10111110100000010011001000100001, 32'b10111110100000010101001010011011, 32'b10111110100000010111001100100000, 32'b10111110100000011001001110110010, 32'b10111110100000011011010001010000, 32'b10111110100000011101010011111010, 32'b10111110100000011111010110110001, 32'b10111110100000100001011001110100, 32'b10111110100000100011011101000011, 32'b10111110100000100101100000011111, 32'b10111110100000100111100100000111, 32'b10111110100000101001100111111100, 32'b10111110100000101011101011111101, 32'b10111110100000101101110000001011, 32'b10111110100000101111110100100101, 32'b10111110100000110001111001001100, 32'b10111110100000110011111110000000, 32'b10111110100000110110000011000000, 32'b10111110100000111000001000001101, 32'b10111110100000111010001101100110, 32'b10111110100000111100010011001100, 32'b10111110100000111110011000111111, 32'b10111110100001000000011110111111, 32'b10111110100001000010100101001011, 32'b10111110100001000100101011100100, 32'b10111110100001000110110010001010, 32'b10111110100001001000111000111101, 32'b10111110100001001010111111111100, 32'b10111110100001001101000111001001, 32'b10111110100001001111001110100010, 32'b10111110100001010001010110001001, 32'b10111110100001010011011101111100, 32'b10111110100001010101100101111100, 32'b10111110100001010111101110001010, 32'b10111110100001011001110110100100, 32'b10111110100001011011111111001100, 32'b10111110100001011110001000000000, 32'b10111110100001100000010001000010, 32'b10111110100001100010011010010001, 32'b10111110100001100100100011101101, 32'b10111110100001100110101101010111, 32'b10111110100001101000110111001101, 32'b10111110100001101011000001010001, 32'b10111110100001101101001011100010, 32'b10111110100001101111010110000000, 32'b10111110100001110001100000101100, 32'b10111110100001110011101011100101, 32'b10111110100001110101110110101100, 32'b10111110100001111000000010000000, 32'b10111110100001111010001101100001, 32'b10111110100001111100011001010000, 32'b10111110100001111110100101001100, 32'b10111110100010000000110001010110, 32'b10111110100010000010111101101110, 32'b10111110100010000101001010010011, 32'b10111110100010000111010111000101, 32'b10111110100010001001100100000101, 32'b10111110100010001011110001010011, 32'b10111110100010001101111110101111, 32'b10111110100010010000001100011000, 32'b10111110100010010010011010001111, 32'b10111110100010010100101000010100, 32'b10111110100010010110110110100111, 32'b10111110100010011001000101000111, 32'b10111110100010011011010011110110, 32'b10111110100010011101100010110010, 32'b10111110100010011111110001111100, 32'b10111110100010100010000001010100, 32'b10111110100010100100010000111010, 32'b10111110100010100110100000101111, 32'b10111110100010101000110000110001, 32'b10111110100010101011000001000001, 32'b10111110100010101101010001011111, 32'b10111110100010101111100010001100, 32'b10111110100010110001110011000110, 32'b10111110100010110100000100001111, 32'b10111110100010110110010101100110, 32'b10111110100010111000100111001011, 32'b10111110100010111010111000111110, 32'b10111110100010111101001011000000, 32'b10111110100010111111011101010000, 32'b10111110100011000001101111101110, 32'b10111110100011000100000010011011, 32'b10111110100011000110010101010110, 32'b10111110100011001000101000100000, 32'b10111110100011001010111011111000, 32'b10111110100011001101001111011110, 32'b10111110100011001111100011010100, 32'b10111110100011010001110111010111, 32'b10111110100011010100001011101001, 32'b10111110100011010110100000001010, 32'b10111110100011011000110100111010, 32'b10111110100011011011001001111000, 32'b10111110100011011101011111000101, 32'b10111110100011011111110100100000, 32'b10111110100011100010001010001011, 32'b10111110100011100100100000000100, 32'b10111110100011100110110110001100, 32'b10111110100011101001001100100011, 32'b10111110100011101011100011001000, 32'b10111110100011101101111001111101, 32'b10111110100011110000010001000001, 32'b10111110100011110010101000010011, 32'b10111110100011110100111111110101, 32'b10111110100011110111010111100101, 32'b10111110100011111001101111100101, 32'b10111110100011111100000111110100, 32'b10111110100011111110100000010010, 32'b10111110100100000000111000111111, 32'b10111110100100000011010001111011, 32'b10111110100100000101101011000111, 32'b10111110100100001000000100100010, 32'b10111110100100001010011110001100, 32'b10111110100100001100111000000101, 32'b10111110100100001111010010001110, 32'b10111110100100010001101100100110, 32'b10111110100100010100000111001110, 32'b10111110100100010110100010000101, 32'b10111110100100011000111101001011, 32'b10111110100100011011011000100001, 32'b10111110100100011101110100000111, 32'b10111110100100100000001111111100, 32'b10111110100100100010101100000001, 32'b10111110100100100101001000010101, 32'b10111110100100100111100100111010, 32'b10111110100100101010000001101101, 32'b10111110100100101100011110110001, 32'b10111110100100101110111100000100, 32'b10111110100100110001011001101000, 32'b10111110100100110011110111011011, 32'b10111110100100110110010101011110, 32'b10111110100100111000110011110000, 32'b10111110100100111011010010010011, 32'b10111110100100111101110001000110, 32'b10111110100101000000010000001001, 32'b10111110100101000010101111011011, 32'b10111110100101000101001110111110, 32'b10111110100101000111101110110001, 32'b10111110100101001010001110110100, 32'b10111110100101001100101111001000, 32'b10111110100101001111001111101011, 32'b10111110100101010001110000011111, 32'b10111110100101010100010001100011, 32'b10111110100101010110110010111000, 32'b10111110100101011001010100011100, 32'b10111110100101011011110110010010, 32'b10111110100101011110011000010111, 32'b10111110100101100000111010101101, 32'b10111110100101100011011101010100, 32'b10111110100101100110000000001011, 32'b10111110100101101000100011010010, 32'b10111110100101101011000110101011, 32'b10111110100101101101101010010011, 32'b10111110100101110000001110001101, 32'b10111110100101110010110010010111, 32'b10111110100101110101010110110010, 32'b10111110100101110111111011011110, 32'b10111110100101111010100000011010, 32'b10111110100101111101000101101000, 32'b10111110100101111111101011000110, 32'b10111110100110000010010000110101, 32'b10111110100110000100110110110101, 32'b10111110100110000111011101000110, 32'b10111110100110001010000011101000, 32'b10111110100110001100101010011100, 32'b10111110100110001111010001100000, 32'b10111110100110010001111000110101, 32'b10111110100110010100100000011100, 32'b10111110100110010111001000010100, 32'b10111110100110011001110000011101, 32'b10111110100110011100011000110111, 32'b10111110100110011111000001100011, 32'b10111110100110100001101010100000, 32'b10111110100110100100010011101110, 32'b10111110100110100110111101001110, 32'b10111110100110101001100110111111, 32'b10111110100110101100010001000010, 32'b10111110100110101110111011010111, 32'b10111110100110110001100101111101, 32'b10111110100110110100010000110100, 32'b10111110100110110110111011111101, 32'b10111110100110111001100111011000, 32'b10111110100110111100010011000101, 32'b10111110100110111110111111000011, 32'b10111110100111000001101011010100, 32'b10111110100111000100010111110110, 32'b10111110100111000111000100101010, 32'b10111110100111001001110001101111, 32'b10111110100111001100011111000111, 32'b10111110100111001111001100110001, 32'b10111110100111010001111010101101, 32'b10111110100111010100101000111011, 32'b10111110100111010111010111011011, 32'b10111110100111011010000110001101, 32'b10111110100111011100110101010010, 32'b10111110100111011111100100101001, 32'b10111110100111100010010100010010, 32'b10111110100111100101000100001101, 32'b10111110100111100111110100011010, 32'b10111110100111101010100100111011, 32'b10111110100111101101010101101101, 32'b10111110100111110000000110110010, 32'b10111110100111110010111000001001, 32'b10111110100111110101101001110011, 32'b10111110100111111000011011110000, 32'b10111110100111111011001101111111, 32'b10111110100111111110000000100001, 32'b10111110101000000000110011010110, 32'b10111110101000000011100110011101, 32'b10111110101000000110011001111000, 32'b10111110101000001001001101100101, 32'b10111110101000001100000001100101, 32'b10111110101000001110110101111000, 32'b10111110101000010001101010011110, 32'b10111110101000010100011111010110, 32'b10111110101000010111010100100010, 32'b10111110101000011010001010000001, 32'b10111110101000011100111111110011, 32'b10111110101000011111110101111001, 32'b10111110101000100010101100010001, 32'b10111110101000100101100010111101, 32'b10111110101000101000011001111100, 32'b10111110101000101011010001001111, 32'b10111110101000101110001000110101, 32'b10111110101000110001000000101110, 32'b10111110101000110011111000111011, 32'b10111110101000110110110001011011, 32'b10111110101000111001101010001111, 32'b10111110101000111100100011010110, 32'b10111110101000111111011100110001, 32'b10111110101001000010010110100000, 32'b10111110101001000101010000100011, 32'b10111110101001001000001010111001, 32'b10111110101001001011000101100011, 32'b10111110101001001110000000100001, 32'b10111110101001010000111011110011, 32'b10111110101001010011110111011001, 32'b10111110101001010110110011010011, 32'b10111110101001011001101111100000, 32'b10111110101001011100101100000010, 32'b10111110101001011111101000111001, 32'b10111110101001100010100110000011, 32'b10111110101001100101100011100001, 32'b10111110101001101000100001010100, 32'b10111110101001101011011111011011, 32'b10111110101001101110011101110111, 32'b10111110101001110001011100100110, 32'b10111110101001110100011011101011, 32'b10111110101001110111011011000100, 32'b10111110101001111010011010110001, 32'b10111110101001111101011010110011, 32'b10111110101010000000011011001001, 32'b10111110101010000011011011110101, 32'b10111110101010000110011100110101, 32'b10111110101010001001011110001001, 32'b10111110101010001100011111110011, 32'b10111110101010001111100001110001, 32'b10111110101010010010100100000101, 32'b10111110101010010101100110101101, 32'b10111110101010011000101001101010, 32'b10111110101010011011101100111100, 32'b10111110101010011110110000100100, 32'b10111110101010100001110100100000, 32'b10111110101010100100111000110010, 32'b10111110101010100111111101011001, 32'b10111110101010101011000010010110, 32'b10111110101010101110000111100111, 32'b10111110101010110001001101001110, 32'b10111110101010110100010011001011, 32'b10111110101010110111011001011101, 32'b10111110101010111010100000000100, 32'b10111110101010111101100111000001, 32'b10111110101011000000101110010100, 32'b10111110101011000011110101111100, 32'b10111110101011000110111101111010, 32'b10111110101011001010000110001110, 32'b10111110101011001101001110111000, 32'b10111110101011010000010111111000, 32'b10111110101011010011100001001101, 32'b10111110101011010110101010111001, 32'b10111110101011011001110100111010, 32'b10111110101011011100111111010010, 32'b10111110101011100000001001111111, 32'b10111110101011100011010101000011, 32'b10111110101011100110100000011101, 32'b10111110101011101001101100001110, 32'b10111110101011101100111000010101, 32'b10111110101011110000000100110010, 32'b10111110101011110011010001100101, 32'b10111110101011110110011110101111, 32'b10111110101011111001101100010000, 32'b10111110101011111100111010000111, 32'b10111110101100000000001000010101, 32'b10111110101100000011010110111001, 32'b10111110101100000110100101110101, 32'b10111110101100001001110101000111, 32'b10111110101100001101000100101111, 32'b10111110101100010000010100101111, 32'b10111110101100010011100101000110, 32'b10111110101100010110110101110100, 32'b10111110101100011010000110111000, 32'b10111110101100011101011000010100, 32'b10111110101100100000101010000111, 32'b10111110101100100011111100010010, 32'b10111110101100100111001110110011, 32'b10111110101100101010100001101100, 32'b10111110101100101101110100111100, 32'b10111110101100110001001000100100, 32'b10111110101100110100011100100011, 32'b10111110101100110111110000111010, 32'b10111110101100111011000101101000, 32'b10111110101100111110011010101110, 32'b10111110101101000001110000001100, 32'b10111110101101000101000110000001, 32'b10111110101101001000011100001110, 32'b10111110101101001011110010110011, 32'b10111110101101001111001001110000, 32'b10111110101101010010100001000101, 32'b10111110101101010101111000110010, 32'b10111110101101011001010000110111, 32'b10111110101101011100101001010101, 32'b10111110101101100000000010001010, 32'b10111110101101100011011011011000, 32'b10111110101101100110110100111110, 32'b10111110101101101010001110111100, 32'b10111110101101101101101001010011, 32'b10111110101101110001000100000011, 32'b10111110101101110100011111001011, 32'b10111110101101110111111010101011, 32'b10111110101101111011010110100100, 32'b10111110101101111110110010110110, 32'b10111110101110000010001111100001, 32'b10111110101110000101101100100100, 32'b10111110101110001001001010000001, 32'b10111110101110001100100111110110, 32'b10111110101110010000000110000100, 32'b10111110101110010011100100101100, 32'b10111110101110010111000011101100, 32'b10111110101110011010100011000110, 32'b10111110101110011110000010111001, 32'b10111110101110100001100011000101, 32'b10111110101110100101000011101011, 32'b10111110101110101000100100101010, 32'b10111110101110101100000110000010, 32'b10111110101110101111100111110101, 32'b10111110101110110011001010000000, 32'b10111110101110110110101100100110, 32'b10111110101110111010001111100101, 32'b10111110101110111101110010111110, 32'b10111110101111000001010110110000, 32'b10111110101111000100111010111101, 32'b10111110101111001000011111100100, 32'b10111110101111001100000100100100, 32'b10111110101111001111101001111111, 32'b10111110101111010011001111110100, 32'b10111110101111010110110110000011, 32'b10111110101111011010011100101100, 32'b10111110101111011110000011110000, 32'b10111110101111100001101011001110, 32'b10111110101111100101010011000111, 32'b10111110101111101000111011011010, 32'b10111110101111101100100100001000, 32'b10111110101111110000001101010000, 32'b10111110101111110011110110110011, 32'b10111110101111110111100000110001, 32'b10111110101111111011001011001010, 32'b10111110101111111110110101111110, 32'b10111110110000000010100001001100, 32'b10111110110000000110001100110110, 32'b10111110110000001001111000111011, 32'b10111110110000001101100101011011, 32'b10111110110000010001010010010110, 32'b10111110110000010100111111101101, 32'b10111110110000011000101101011111, 32'b10111110110000011100011011101100, 32'b10111110110000100000001010010101, 32'b10111110110000100011111001011001, 32'b10111110110000100111101000111001, 32'b10111110110000101011011000110101, 32'b10111110110000101111001001001101, 32'b10111110110000110010111010000000, 32'b10111110110000110110101011001111, 32'b10111110110000111010011100111010, 32'b10111110110000111110001111000010, 32'b10111110110001000010000001100101, 32'b10111110110001000101110100100101, 32'b10111110110001001001101000000000, 32'b10111110110001001101011011111000, 32'b10111110110001010001010000001101, 32'b10111110110001010101000100111110, 32'b10111110110001011000111010001011, 32'b10111110110001011100101111110101, 32'b10111110110001100000100101111100, 32'b10111110110001100100011100011111, 32'b10111110110001101000010011100000, 32'b10111110110001101100001010111101, 32'b10111110110001110000000010110111, 32'b10111110110001110011111011001110, 32'b10111110110001110111110100000010, 32'b10111110110001111011101101010011, 32'b10111110110001111111100111000001, 32'b10111110110010000011100001001101, 32'b10111110110010000111011011110110, 32'b10111110110010001011010110111101, 32'b10111110110010001111010010100001, 32'b10111110110010010011001110100010, 32'b10111110110010010111001011000010, 32'b10111110110010011011000111111111, 32'b10111110110010011111000101011001, 32'b10111110110010100011000011010010, 32'b10111110110010100111000001101001, 32'b10111110110010101011000000011101, 32'b10111110110010101110111111110000, 32'b10111110110010110010111111100001, 32'b10111110110010110110111111110000, 32'b10111110110010111011000000011101, 32'b10111110110010111111000001101001, 32'b10111110110011000011000011010011, 32'b10111110110011000111000101011100, 32'b10111110110011001011001000000100, 32'b10111110110011001111001011001010, 32'b10111110110011010011001110101110, 32'b10111110110011010111010010110010, 32'b10111110110011011011010111010101, 32'b10111110110011011111011100010110, 32'b10111110110011100011100001110111, 32'b10111110110011100111100111110111, 32'b10111110110011101011101110010110, 32'b10111110110011101111110101010100, 32'b10111110110011110011111100110010, 32'b10111110110011111000000100101111, 32'b10111110110011111100001101001100, 32'b10111110110100000000010110001000, 32'b10111110110100000100011111100100, 32'b10111110110100001000101001100000, 32'b10111110110100001100110011111100, 32'b10111110110100010000111110110111, 32'b10111110110100010101001010010011, 32'b10111110110100011001010110001111, 32'b10111110110100011101100010101011, 32'b10111110110100100001101111100111, 32'b10111110110100100101111101000011, 32'b10111110110100101010001011000000, 32'b10111110110100101110011001011101, 32'b10111110110100110010101000011011, 32'b10111110110100110110110111111010, 32'b10111110110100111011000111111001, 32'b10111110110100111111011000011010, 32'b10111110110101000011101001011011, 32'b10111110110101000111111010111101, 32'b10111110110101001100001101000000, 32'b10111110110101010000011111100100, 32'b10111110110101010100110010101010, 32'b10111110110101011001000110010001, 32'b10111110110101011101011010011001, 32'b10111110110101100001101111000011, 32'b10111110110101100110000100001110, 32'b10111110110101101010011001111011, 32'b10111110110101101110110000001010, 32'b10111110110101110011000110111010, 32'b10111110110101110111011110001101, 32'b10111110110101111011110110000001, 32'b10111110110110000000001110011000, 32'b10111110110110000100100111010001, 32'b10111110110110001001000000101100, 32'b10111110110110001101011010101001, 32'b10111110110110010001110101001001, 32'b10111110110110010110010000001011, 32'b10111110110110011010101011110000, 32'b10111110110110011111000111111000, 32'b10111110110110100011100100100010, 32'b10111110110110101000000001101111, 32'b10111110110110101100011111100000, 32'b10111110110110110000111101110011, 32'b10111110110110110101011100101010, 32'b10111110110110111001111100000011, 32'b10111110110110111110011100000000, 32'b10111110110111000010111100100001, 32'b10111110110111000111011101100101, 32'b10111110110111001011111111001100, 32'b10111110110111010000100001011000, 32'b10111110110111010101000100000111, 32'b10111110110111011001100111011010, 32'b10111110110111011110001011010000, 32'b10111110110111100010101111101011, 32'b10111110110111100111010100101011, 32'b10111110110111101011111010001110, 32'b10111110110111110000100000010110, 32'b10111110110111110101000111000010, 32'b10111110110111111001101110010010, 32'b10111110110111111110010110001000, 32'b10111110111000000010111110100010, 32'b10111110111000000111100111100000, 32'b10111110111000001100010001000100, 32'b10111110111000010000111011001101, 32'b10111110111000010101100101111011, 32'b10111110111000011010010001001110, 32'b10111110111000011110111101000110, 32'b10111110111000100011101001100100, 32'b10111110111000101000010110100111, 32'b10111110111000101101000100010000, 32'b10111110111000110001110010011110, 32'b10111110111000110110100001010010, 32'b10111110111000111011010000101100, 32'b10111110111001000000000000101100, 32'b10111110111001000100110001010010, 32'b10111110111001001001100010011111, 32'b10111110111001001110010100010001, 32'b10111110111001010011000110101010, 32'b10111110111001010111111001101010, 32'b10111110111001011100101101010000, 32'b10111110111001100001100001011100, 32'b10111110111001100110010110010000, 32'b10111110111001101011001011101010, 32'b10111110111001110000000001101011, 32'b10111110111001110100111000010100, 32'b10111110111001111001101111100011, 32'b10111110111001111110100111011010, 32'b10111110111010000011011111111001, 32'b10111110111010001000011000111110, 32'b10111110111010001101010010101100, 32'b10111110111010010010001101000001, 32'b10111110111010010111000111111110, 32'b10111110111010011100000011100010, 32'b10111110111010100000111111101111, 32'b10111110111010100101111100100100, 32'b10111110111010101010111010000001, 32'b10111110111010101111111000000111, 32'b10111110111010110100110110110101, 32'b10111110111010111001110110001011, 32'b10111110111010111110110110001011, 32'b10111110111011000011110110110010, 32'b10111110111011001000111000000011, 32'b10111110111011001101111001111101, 32'b10111110111011010010111100100000, 32'b10111110111011010111111111101100, 32'b10111110111011011101000011100001, 32'b10111110111011100010001000000000, 32'b10111110111011100111001101001001, 32'b10111110111011101100010010111011, 32'b10111110111011110001011001010110, 32'b10111110111011110110100000011100, 32'b10111110111011111011101000001100, 32'b10111110111100000000110000100101, 32'b10111110111100000101111001101001, 32'b10111110111100001011000011010111, 32'b10111110111100010000001101110000, 32'b10111110111100010101011000110011, 32'b10111110111100011010100100100001, 32'b10111110111100011111110000111010, 32'b10111110111100100100111101111101, 32'b10111110111100101010001011101100, 32'b10111110111100101111011010000110, 32'b10111110111100110100101001001010, 32'b10111110111100111001111000111011, 32'b10111110111100111111001001010110, 32'b10111110111101000100011010011110, 32'b10111110111101001001101100010001, 32'b10111110111101001110111110101111, 32'b10111110111101010100010001111010, 32'b10111110111101011001100101110001, 32'b10111110111101011110111010010100, 32'b10111110111101100100001111100011, 32'b10111110111101101001100101011111, 32'b10111110111101101110111100000111, 32'b10111110111101110100010011011100, 32'b10111110111101111001101011011110, 32'b10111110111101111111000100001100, 32'b10111110111110000100011101101000, 32'b10111110111110001001110111110001, 32'b10111110111110001111010010100111, 32'b10111110111110010100101110001010, 32'b10111110111110011010001010011011, 32'b10111110111110011111100111011010, 32'b10111110111110100101000101000110, 32'b10111110111110101010100011100000, 32'b10111110111110110000000010101001, 32'b10111110111110110101100010011111, 32'b10111110111110111011000011000100, 32'b10111110111111000000100100010111, 32'b10111110111111000110000110011001, 32'b10111110111111001011101001001001, 32'b10111110111111010001001100101000, 32'b10111110111111010110110000110110, 32'b10111110111111011100010101110011, 32'b10111110111111100001111011011111, 32'b10111110111111100111100001111010, 32'b10111110111111101101001001000101, 32'b10111110111111110010110001000000, 32'b10111110111111111000011001101010, 32'b10111110111111111110000011000100, 32'b10111111000000000001110110100111, 32'b10111111000000000100101100000100, 32'b10111111000000000111100001111001, 32'b10111111000000001010011000000110, 32'b10111111000000001101001110101100, 32'b10111111000000010000000101101010, 32'b10111111000000010010111101000000, 32'b10111111000000010101110100101111, 32'b10111111000000011000101100110110, 32'b10111111000000011011100101010101, 32'b10111111000000011110011110001110, 32'b10111111000000100001010111011111, 32'b10111111000000100100010001001001, 32'b10111111000000100111001011001100, 32'b10111111000000101010000101100111, 32'b10111111000000101101000000011100, 32'b10111111000000101111111011101010, 32'b10111111000000110010110111010001, 32'b10111111000000110101110011010001, 32'b10111111000000111000101111101010, 32'b10111111000000111011101100011101, 32'b10111111000000111110101001101001, 32'b10111111000001000001100111001111, 32'b10111111000001000100100101001110, 32'b10111111000001000111100011100111, 32'b10111111000001001010100010011001, 32'b10111111000001001101100001100110, 32'b10111111000001010000100001001100, 32'b10111111000001010011100001001100, 32'b10111111000001010110100001100110, 32'b10111111000001011001100010011010, 32'b10111111000001011100100011101001, 32'b10111111000001011111100101010001, 32'b10111111000001100010100111010100, 32'b10111111000001100101101001110001, 32'b10111111000001101000101100101001, 32'b10111111000001101011101111111011, 32'b10111111000001101110110011101000, 32'b10111111000001110001110111101111, 32'b10111111000001110100111100010001, 32'b10111111000001111000000001001110, 32'b10111111000001111011000110100110, 32'b10111111000001111110001100011001, 32'b10111111000010000001010010100111, 32'b10111111000010000100011001010000, 32'b10111111000010000111100000010100, 32'b10111111000010001010100111110100, 32'b10111111000010001101101111101111, 32'b10111111000010010000111000000101, 32'b10111111000010010100000000110111, 32'b10111111000010010111001010000100, 32'b10111111000010011010010011101101, 32'b10111111000010011101011101110010, 32'b10111111000010100000101000010011, 32'b10111111000010100011110011001111, 32'b10111111000010100110111110101000, 32'b10111111000010101010001010011100, 32'b10111111000010101101010110101101, 32'b10111111000010110000100011011010, 32'b10111111000010110011110000100100, 32'b10111111000010110110111110001001, 32'b10111111000010111010001100001100, 32'b10111111000010111101011010101010, 32'b10111111000011000000101001100110, 32'b10111111000011000011111000111110, 32'b10111111000011000111001000110011, 32'b10111111000011001010011001000101, 32'b10111111000011001101101001110100, 32'b10111111000011010000111011000000, 32'b10111111000011010100001100101001, 32'b10111111000011010111011110101111, 32'b10111111000011011010110001010011, 32'b10111111000011011110000100010100, 32'b10111111000011100001010111110010, 32'b10111111000011100100101011101110, 32'b10111111000011101000000000001000, 32'b10111111000011101011010100111111, 32'b10111111000011101110101010010101, 32'b10111111000011110010000000001000, 32'b10111111000011110101010110011001, 32'b10111111000011111000101101001000, 32'b10111111000011111100000100010110, 32'b10111111000011111111011100000010, 32'b10111111000100000010110100001100, 32'b10111111000100000110001100110100, 32'b10111111000100001001100101111100, 32'b10111111000100001100111111100001, 32'b10111111000100010000011001100110, 32'b10111111000100010011110100001001, 32'b10111111000100010111001111001011, 32'b10111111000100011010101010101100, 32'b10111111000100011110000110101101, 32'b10111111000100100001100011001100, 32'b10111111000100100101000000001011, 32'b10111111000100101000011101101001, 32'b10111111000100101011111011100110, 32'b10111111000100101111011010000011, 32'b10111111000100110010111001000000, 32'b10111111000100110110011000011100, 32'b10111111000100111001111000011001, 32'b10111111000100111101011000110101, 32'b10111111000101000000111001110001, 32'b10111111000101000100011011001101, 32'b10111111000101000111111101001010, 32'b10111111000101001011011111100111, 32'b10111111000101001111000010100100, 32'b10111111000101010010100110000010, 32'b10111111000101010110001010000000, 32'b10111111000101011001101110011111, 32'b10111111000101011101010011011111, 32'b10111111000101100000111000111111, 32'b10111111000101100100011111000001, 32'b10111111000101101000000101100100, 32'b10111111000101101011101100100111, 32'b10111111000101101111010100001101, 32'b10111111000101110010111100010011, 32'b10111111000101110110100100111011, 32'b10111111000101111010001110000101, 32'b10111111000101111101110111110000, 32'b10111111000110000001100001111101, 32'b10111111000110000101001100101100, 32'b10111111000110001000110111111101, 32'b10111111000110001100100011110000, 32'b10111111000110010000010000000101, 32'b10111111000110010011111100111101, 32'b10111111000110010111101010010111, 32'b10111111000110011011011000010011, 32'b10111111000110011111000110110010, 32'b10111111000110100010110101110100, 32'b10111111000110100110100101011001, 32'b10111111000110101010010101100000, 32'b10111111000110101110000110001011, 32'b10111111000110110001110111011001, 32'b10111111000110110101101001001001, 32'b10111111000110111001011011011110, 32'b10111111000110111101001110010110, 32'b10111111000111000001000001110001, 32'b10111111000111000100110101110000, 32'b10111111000111001000101010010011, 32'b10111111000111001100011111011001, 32'b10111111000111010000010101000100, 32'b10111111000111010100001011010011, 32'b10111111000111011000000010000110, 32'b10111111000111011011111001011101, 32'b10111111000111011111110001011001, 32'b10111111000111100011101001111001, 32'b10111111000111100111100010111110, 32'b10111111000111101011011100101000, 32'b10111111000111101111010110110111, 32'b10111111000111110011010001101011, 32'b10111111000111110111001101000100, 32'b10111111000111111011001001000010, 32'b10111111000111111111000101100101, 32'b10111111001000000011000010101110, 32'b10111111001000000111000000011101, 32'b10111111001000001010111110110001, 32'b10111111001000001110111101101011, 32'b10111111001000010010111101001011, 32'b10111111001000010110111101010001, 32'b10111111001000011010111101111110, 32'b10111111001000011110111111010000, 32'b10111111001000100011000001001001, 32'b10111111001000100111000011101001, 32'b10111111001000101011000110101111, 32'b10111111001000101111001010011100, 32'b10111111001000110011001110101111, 32'b10111111001000110111010011101010, 32'b10111111001000111011011001001100, 32'b10111111001000111111011111010101, 32'b10111111001001000011100110000110, 32'b10111111001001000111101101011110, 32'b10111111001001001011110101011110, 32'b10111111001001001111111110000101, 32'b10111111001001010100000111010101, 32'b10111111001001011000010001001100, 32'b10111111001001011100011011101100, 32'b10111111001001100000100110110011, 32'b10111111001001100100110010100100, 32'b10111111001001101000111110111100, 32'b10111111001001101101001011111110, 32'b10111111001001110001011001101000, 32'b10111111001001110101100111111011, 32'b10111111001001111001110110110111, 32'b10111111001001111110000110011100, 32'b10111111001010000010010110101010, 32'b10111111001010000110100111100010, 32'b10111111001010001010111001000011, 32'b10111111001010001111001011001111, 32'b10111111001010010011011110000011, 32'b10111111001010010111110001100010, 32'b10111111001010011100000101101011, 32'b10111111001010100000011010011110, 32'b10111111001010100100101111111100, 32'b10111111001010101001000110000100, 32'b10111111001010101101011100110110, 32'b10111111001010110001110100010100, 32'b10111111001010110110001100011100, 32'b10111111001010111010100101001111, 32'b10111111001010111110111110101101, 32'b10111111001011000011011000110111, 32'b10111111001011000111110011101100, 32'b10111111001011001100001111001101, 32'b10111111001011010000101011011010, 32'b10111111001011010101001000010010, 32'b10111111001011011001100101110110, 32'b10111111001011011110000100000111, 32'b10111111001011100010100011000011, 32'b10111111001011100111000010101101, 32'b10111111001011101011100011000010, 32'b10111111001011110000000100000101, 32'b10111111001011110100100101110100, 32'b10111111001011111001001000010001, 32'b10111111001011111101101011011010, 32'b10111111001100000010001111010001, 32'b10111111001100000110110011110101, 32'b10111111001100001011011001000111, 32'b10111111001100001111111111000111, 32'b10111111001100010100100101110100, 32'b10111111001100011001001101010000, 32'b10111111001100011101110101011001, 32'b10111111001100100010011110010001, 32'b10111111001100100111000111111000, 32'b10111111001100101011110010001101, 32'b10111111001100110000011101010001, 32'b10111111001100110101001001000100, 32'b10111111001100111001110101100110, 32'b10111111001100111110100010110111, 32'b10111111001101000011010000111000, 32'b10111111001101000111111111101000, 32'b10111111001101001100101111001000, 32'b10111111001101010001011111011000, 32'b10111111001101010110010000011000, 32'b10111111001101011011000010001000, 32'b10111111001101011111110100101001, 32'b10111111001101100100100111111010, 32'b10111111001101101001011011111100, 32'b10111111001101101110010000101110, 32'b10111111001101110011000110010010, 32'b10111111001101110111111100100110, 32'b10111111001101111100110011101100, 32'b10111111001110000001101011100100, 32'b10111111001110000110100100001101, 32'b10111111001110001011011101101000, 32'b10111111001110010000010111110101, 32'b10111111001110010101010010110100, 32'b10111111001110011010001110100101, 32'b10111111001110011111001011001001, 32'b10111111001110100100001000100000, 32'b10111111001110101001000110101001, 32'b10111111001110101110000101100101, 32'b10111111001110110011000101010101, 32'b10111111001110111000000101111000, 32'b10111111001110111101000111001110, 32'b10111111001111000010001001011000, 32'b10111111001111000111001100010110, 32'b10111111001111001100010000001000, 32'b10111111001111010001010100101110, 32'b10111111001111010110011010001000, 32'b10111111001111011011100000010111, 32'b10111111001111100000100111011011, 32'b10111111001111100101101111010011, 32'b10111111001111101010111000000001, 32'b10111111001111110000000001100100, 32'b10111111001111110101001011111100, 32'b10111111001111111010010111001010, 32'b10111111001111111111100011001110, 32'b10111111010000000100110000001000, 32'b10111111010000001001111101111000, 32'b10111111010000001111001100011110, 32'b10111111010000010100011011111011, 32'b10111111010000011001101100001111, 32'b10111111010000011110111101011001, 32'b10111111010000100100001111011011, 32'b10111111010000101001100010010100, 32'b10111111010000101110110110000100, 32'b10111111010000110100001010101100, 32'b10111111010000111001100000001100, 32'b10111111010000111110110110100100, 32'b10111111010001000100001101110100, 32'b10111111010001001001100101111100, 32'b10111111010001001110111110111101, 32'b10111111010001010100011000110111, 32'b10111111010001011001110011101010, 32'b10111111010001011111001111010111, 32'b10111111010001100100101011111100, 32'b10111111010001101010001001011011, 32'b10111111010001101111100111110100, 32'b10111111010001110101000111000111, 32'b10111111010001111010100111010100, 32'b10111111010010000000001000011100, 32'b10111111010010000101101010011110, 32'b10111111010010001011001101011011, 32'b10111111010010010000110001010011, 32'b10111111010010010110010110000110, 32'b10111111010010011011111011110101, 32'b10111111010010100001100010011111, 32'b10111111010010100111001010000101, 32'b10111111010010101100110010100111, 32'b10111111010010110010011100000101, 32'b10111111010010111000000110100000, 32'b10111111010010111101110001110111, 32'b10111111010011000011011110001100, 32'b10111111010011001001001011011101, 32'b10111111010011001110111001101100, 32'b10111111010011010100101000111000, 32'b10111111010011011010011001000010, 32'b10111111010011100000001010001010, 32'b10111111010011100101111100010000, 32'b10111111010011101011101111010101, 32'b10111111010011110001100011011000, 32'b10111111010011110111011000011010, 32'b10111111010011111101001110011010, 32'b10111111010100000011000101011011, 32'b10111111010100001000111101011010, 32'b10111111010100001110110110011010, 32'b10111111010100010100110000011001, 32'b10111111010100011010101011011001, 32'b10111111010100100000100111011001, 32'b10111111010100100110100100011001, 32'b10111111010100101100100010011011, 32'b10111111010100110010100001011101, 32'b10111111010100111000100001100001, 32'b10111111010100111110100010100110, 32'b10111111010101000100100100101101, 32'b10111111010101001010100111110111, 32'b10111111010101010000101100000010, 32'b10111111010101010110110001010000, 32'b10111111010101011100110111100000, 32'b10111111010101100010111110110100, 32'b10111111010101101001000111001011, 32'b10111111010101101111010000100101, 32'b10111111010101110101011011000011, 32'b10111111010101111011100110100101, 32'b10111111010110000001110011001011, 32'b10111111010110001000000000110101, 32'b10111111010110001110001111100100, 32'b10111111010110010100011111011000, 32'b10111111010110011010110000010001, 32'b10111111010110100001000010010000, 32'b10111111010110100111010101010100, 32'b10111111010110101101101001011110, 32'b10111111010110110011111110101110, 32'b10111111010110111010010101000101, 32'b10111111010111000000101100100010, 32'b10111111010111000111000101000111, 32'b10111111010111001101011110110010, 32'b10111111010111010011111001100101, 32'b10111111010111011010010101011111, 32'b10111111010111100000110010100010, 32'b10111111010111100111010000101101, 32'b10111111010111101101110000000000, 32'b10111111010111110100010000011100, 32'b10111111010111111010110010000001, 32'b10111111011000000001010100110000, 32'b10111111011000000111111000100111, 32'b10111111011000001110011101101001, 32'b10111111011000010101000011110101, 32'b10111111011000011011101011001011, 32'b10111111011000100010010011101100, 32'b10111111011000101000111101011000, 32'b10111111011000101111101000001111, 32'b10111111011000110110010100010001, 32'b10111111011000111101000001011111, 32'b10111111011001000011101111111001, 32'b10111111011001001010011111100000, 32'b10111111011001010001010000010011, 32'b10111111011001011000000010010011, 32'b10111111011001011110110101100000, 32'b10111111011001100101101001111010, 32'b10111111011001101100011111100010, 32'b10111111011001110011010110011001, 32'b10111111011001111010001110011101, 32'b10111111011010000001000111110000, 32'b10111111011010001000000010010011, 32'b10111111011010001110111110000100, 32'b10111111011010010101111011000100, 32'b10111111011010011100111001010101, 32'b10111111011010100011111000110110, 32'b10111111011010101010111001100111, 32'b10111111011010110001111011101000, 32'b10111111011010111000111110111011, 32'b10111111011011000000000011011111, 32'b10111111011011000111001001010100, 32'b10111111011011001110010000011011, 32'b10111111011011010101011000110101, 32'b10111111011011011100100010100001, 32'b10111111011011100011101101100000, 32'b10111111011011101010111001110010, 32'b10111111011011110010000111011000, 32'b10111111011011111001010110010001, 32'b10111111011100000000100110011110, 32'b10111111011100000111111000000000, 32'b10111111011100001111001010110110, 32'b10111111011100010110011111000010, 32'b10111111011100011101110100100011, 32'b10111111011100100101001011011001, 32'b10111111011100101100100011100110, 32'b10111111011100110011111101001001, 32'b10111111011100111011011000000011, 32'b10111111011101000010110100010011, 32'b10111111011101001010010001111011, 32'b10111111011101010001110000111011, 32'b10111111011101011001010001010010, 32'b10111111011101100000110011000010, 32'b10111111011101101000010110001011, 32'b10111111011101101111111010101101, 32'b10111111011101110111100000101000, 32'b10111111011101111111000111111101, 32'b10111111011110000110110000101011, 32'b10111111011110001110011010110101, 32'b10111111011110010110000110011001, 32'b10111111011110011101110011011000, 32'b10111111011110100101100001110010, 32'b10111111011110101101010001101000, 32'b10111111011110110101000010111011, 32'b10111111011110111100110101101010, 32'b10111111011111000100101001110110, 32'b10111111011111001100011111011111, 32'b10111111011111010100010110100110, 32'b10111111011111011100001111001010, 32'b10111111011111100100001001001101, 32'b10111111011111101100000100101111, 32'b10111111011111110100000001110000, 32'b10111111011111111100000000010000};


    assign b_table = '{32'b00111111100000000000100000000001, 32'b00111111100000000001100000000101, 32'b00111111100000000010100000001101, 32'b00111111100000000011100000011001, 32'b00111111100000000100100000101001, 32'b00111111100000000101100000111101, 32'b00111111100000000110100001010101, 32'b00111111100000000111100001110001, 32'b00111111100000001000100010010001, 32'b00111111100000001001100010110110, 32'b00111111100000001010100011011110, 32'b00111111100000001011100100001010, 32'b00111111100000001100100100111011, 32'b00111111100000001101100101101111, 32'b00111111100000001110100110101000, 32'b00111111100000001111100111100101, 32'b00111111100000010000101000100101, 32'b00111111100000010001101001101010, 32'b00111111100000010010101010110011, 32'b00111111100000010011101100000000, 32'b00111111100000010100101101010001, 32'b00111111100000010101101110100111, 32'b00111111100000010110110000000000, 32'b00111111100000010111110001011110, 32'b00111111100000011000110010111111, 32'b00111111100000011001110100100101, 32'b00111111100000011010110110001111, 32'b00111111100000011011110111111101, 32'b00111111100000011100111001110000, 32'b00111111100000011101111011100110, 32'b00111111100000011110111101100001, 32'b00111111100000011111111111100000, 32'b00111111100000100001000001100011, 32'b00111111100000100010000011101010, 32'b00111111100000100011000101110110, 32'b00111111100000100100001000000101, 32'b00111111100000100101001010011001, 32'b00111111100000100110001100110001, 32'b00111111100000100111001111001110, 32'b00111111100000101000010001101110, 32'b00111111100000101001010100010011, 32'b00111111100000101010010110111100, 32'b00111111100000101011011001101001, 32'b00111111100000101100011100011011, 32'b00111111100000101101011111010001, 32'b00111111100000101110100010001011, 32'b00111111100000101111100101001001, 32'b00111111100000110000101000001100, 32'b00111111100000110001101011010011, 32'b00111111100000110010101110011110, 32'b00111111100000110011110001101110, 32'b00111111100000110100110101000010, 32'b00111111100000110101111000011010, 32'b00111111100000110110111011110110, 32'b00111111100000110111111111010111, 32'b00111111100000111001000010111101, 32'b00111111100000111010000110100110, 32'b00111111100000111011001010010100, 32'b00111111100000111100001110000110, 32'b00111111100000111101010001111101, 32'b00111111100000111110010101111000, 32'b00111111100000111111011001110111, 32'b00111111100001000000011101111011, 32'b00111111100001000001100010000011, 32'b00111111100001000010100110001111, 32'b00111111100001000011101010100000, 32'b00111111100001000100101110110110, 32'b00111111100001000101110011001111, 32'b00111111100001000110110111101110, 32'b00111111100001000111111100010000, 32'b00111111100001001001000000110111, 32'b00111111100001001010000101100011, 32'b00111111100001001011001010010011, 32'b00111111100001001100001111000111, 32'b00111111100001001101010100000000, 32'b00111111100001001110011000111101, 32'b00111111100001001111011101111111, 32'b00111111100001010000100011000101, 32'b00111111100001010001101000010000, 32'b00111111100001010010101101011111, 32'b00111111100001010011110010110011, 32'b00111111100001010100111000001011, 32'b00111111100001010101111101101000, 32'b00111111100001010111000011001010, 32'b00111111100001011000001000101111, 32'b00111111100001011001001110011010, 32'b00111111100001011010010100001001, 32'b00111111100001011011011001111100, 32'b00111111100001011100011111110100, 32'b00111111100001011101100101110001, 32'b00111111100001011110101011110010, 32'b00111111100001011111110001111000, 32'b00111111100001100000111000000010, 32'b00111111100001100001111110010001, 32'b00111111100001100011000100100101, 32'b00111111100001100100001010111101, 32'b00111111100001100101010001011010, 32'b00111111100001100110010111111011, 32'b00111111100001100111011110100001, 32'b00111111100001101000100101001100, 32'b00111111100001101001101011111011, 32'b00111111100001101010110010101111, 32'b00111111100001101011111001101000, 32'b00111111100001101101000000100101, 32'b00111111100001101110000111100111, 32'b00111111100001101111001110101110, 32'b00111111100001110000010101111001, 32'b00111111100001110001011101001001, 32'b00111111100001110010100100011110, 32'b00111111100001110011101011111000, 32'b00111111100001110100110011010110, 32'b00111111100001110101111010111001, 32'b00111111100001110111000010100000, 32'b00111111100001111000001010001101, 32'b00111111100001111001010001111110, 32'b00111111100001111010011001110100, 32'b00111111100001111011100001101110, 32'b00111111100001111100101001101110, 32'b00111111100001111101110001110010, 32'b00111111100001111110111001111011, 32'b00111111100010000000000010001000, 32'b00111111100010000001001010011011, 32'b00111111100010000010010010110010, 32'b00111111100010000011011011001111, 32'b00111111100010000100100011101111, 32'b00111111100010000101101100010101, 32'b00111111100010000110110101000000, 32'b00111111100010000111111101101111, 32'b00111111100010001001000110100100, 32'b00111111100010001010001111011101, 32'b00111111100010001011011000011011, 32'b00111111100010001100100001011110, 32'b00111111100010001101101010100110, 32'b00111111100010001110110011110010, 32'b00111111100010001111111101000100, 32'b00111111100010010001000110011011, 32'b00111111100010010010001111110110, 32'b00111111100010010011011001010110, 32'b00111111100010010100100010111100, 32'b00111111100010010101101100100110, 32'b00111111100010010110110110010101, 32'b00111111100010011000000000001001, 32'b00111111100010011001001010000010, 32'b00111111100010011010010100000000, 32'b00111111100010011011011110000011, 32'b00111111100010011100101000001011, 32'b00111111100010011101110010011000, 32'b00111111100010011110111100101010, 32'b00111111100010100000000111000001, 32'b00111111100010100001010001011101, 32'b00111111100010100010011011111110, 32'b00111111100010100011100110100100, 32'b00111111100010100100110001001111, 32'b00111111100010100101111011111111, 32'b00111111100010100111000110110100, 32'b00111111100010101000010001101111, 32'b00111111100010101001011100101110, 32'b00111111100010101010100111110010, 32'b00111111100010101011110010111100, 32'b00111111100010101100111110001010, 32'b00111111100010101110001001011110, 32'b00111111100010101111010100110111, 32'b00111111100010110000100000010101, 32'b00111111100010110001101011111000, 32'b00111111100010110010110111100000, 32'b00111111100010110100000011001101, 32'b00111111100010110101001110111111, 32'b00111111100010110110011010110111, 32'b00111111100010110111100110110100, 32'b00111111100010111000110010110110, 32'b00111111100010111001111110111101, 32'b00111111100010111011001011001001, 32'b00111111100010111100010111011011, 32'b00111111100010111101100011110001, 32'b00111111100010111110110000001101, 32'b00111111100010111111111100101110, 32'b00111111100011000001001001010101, 32'b00111111100011000010010110000001, 32'b00111111100011000011100010110001, 32'b00111111100011000100101111101000, 32'b00111111100011000101111100100011, 32'b00111111100011000111001001100100, 32'b00111111100011001000010110101010, 32'b00111111100011001001100011110101, 32'b00111111100011001010110001000101, 32'b00111111100011001011111110011011, 32'b00111111100011001101001011110111, 32'b00111111100011001110011001010111, 32'b00111111100011001111100110111101, 32'b00111111100011010000110100101000, 32'b00111111100011010010000010011001, 32'b00111111100011010011010000001111, 32'b00111111100011010100011110001010, 32'b00111111100011010101101100001011, 32'b00111111100011010110111010010001, 32'b00111111100011011000001000011100, 32'b00111111100011011001010110101101, 32'b00111111100011011010100101000011, 32'b00111111100011011011110011011111, 32'b00111111100011011101000010000000, 32'b00111111100011011110010000100110, 32'b00111111100011011111011111010010, 32'b00111111100011100000101110000100, 32'b00111111100011100001111100111011, 32'b00111111100011100011001011110111, 32'b00111111100011100100011010111001, 32'b00111111100011100101101010000001, 32'b00111111100011100110111001001101, 32'b00111111100011101000001000100000, 32'b00111111100011101001010111111000, 32'b00111111100011101010100111010101, 32'b00111111100011101011110110111000, 32'b00111111100011101101000110100001, 32'b00111111100011101110010110001111, 32'b00111111100011101111100110000010, 32'b00111111100011110000110101111100, 32'b00111111100011110010000101111010, 32'b00111111100011110011010101111111, 32'b00111111100011110100100110001001, 32'b00111111100011110101110110011001, 32'b00111111100011110111000110101110, 32'b00111111100011111000010111001001, 32'b00111111100011111001100111101001, 32'b00111111100011111010111000001111, 32'b00111111100011111100001000111011, 32'b00111111100011111101011001101101, 32'b00111111100011111110101010100100, 32'b00111111100011111111111011100001, 32'b00111111100100000001001100100011, 32'b00111111100100000010011101101011, 32'b00111111100100000011101110111001, 32'b00111111100100000101000000001101, 32'b00111111100100000110010001100110, 32'b00111111100100000111100011000101, 32'b00111111100100001000110100101010, 32'b00111111100100001010000110010101, 32'b00111111100100001011011000000101, 32'b00111111100100001100101001111100, 32'b00111111100100001101111011111000, 32'b00111111100100001111001101111010, 32'b00111111100100010000100000000001, 32'b00111111100100010001110010001111, 32'b00111111100100010011000100100010, 32'b00111111100100010100010110111011, 32'b00111111100100010101101001011010, 32'b00111111100100010110111011111111, 32'b00111111100100011000001110101001, 32'b00111111100100011001100001011010, 32'b00111111100100011010110100010000, 32'b00111111100100011100000111001101, 32'b00111111100100011101011010001111, 32'b00111111100100011110101101010111, 32'b00111111100100100000000000100101, 32'b00111111100100100001010011111001, 32'b00111111100100100010100111010011, 32'b00111111100100100011111010110011, 32'b00111111100100100101001110011001, 32'b00111111100100100110100010000101, 32'b00111111100100100111110101110111, 32'b00111111100100101001001001101110, 32'b00111111100100101010011101101100, 32'b00111111100100101011110001110000, 32'b00111111100100101101000101111010, 32'b00111111100100101110011010001010, 32'b00111111100100101111101110100000, 32'b00111111100100110001000010111100, 32'b00111111100100110010010111011110, 32'b00111111100100110011101100000110, 32'b00111111100100110101000000110100, 32'b00111111100100110110010101101001, 32'b00111111100100110111101010100011, 32'b00111111100100111000111111100100, 32'b00111111100100111010010100101010, 32'b00111111100100111011101001110111, 32'b00111111100100111100111111001010, 32'b00111111100100111110010100100011, 32'b00111111100100111111101010000011, 32'b00111111100101000000111111101000, 32'b00111111100101000010010101010100, 32'b00111111100101000011101011000110, 32'b00111111100101000101000000111110, 32'b00111111100101000110010110111100, 32'b00111111100101000111101101000001, 32'b00111111100101001001000011001100, 32'b00111111100101001010011001011101, 32'b00111111100101001011101111110100, 32'b00111111100101001101000110010010, 32'b00111111100101001110011100110110, 32'b00111111100101001111110011100000, 32'b00111111100101010001001010010000, 32'b00111111100101010010100001000111, 32'b00111111100101010011111000000100, 32'b00111111100101010101001111001000, 32'b00111111100101010110100110010010, 32'b00111111100101010111111101100010, 32'b00111111100101011001010100111000, 32'b00111111100101011010101100010101, 32'b00111111100101011100000011111001, 32'b00111111100101011101011011100010, 32'b00111111100101011110110011010011, 32'b00111111100101100000001011001001, 32'b00111111100101100001100011000110, 32'b00111111100101100010111011001010, 32'b00111111100101100100010011010100, 32'b00111111100101100101101011100100, 32'b00111111100101100111000011111011, 32'b00111111100101101000011100011000, 32'b00111111100101101001110100111100, 32'b00111111100101101011001101100111, 32'b00111111100101101100100110011000, 32'b00111111100101101101111111001111, 32'b00111111100101101111011000001101, 32'b00111111100101110000110001010010, 32'b00111111100101110010001010011101, 32'b00111111100101110011100011101111, 32'b00111111100101110100111101000111, 32'b00111111100101110110010110100110, 32'b00111111100101110111110000001100, 32'b00111111100101111001001001111000, 32'b00111111100101111010100011101011, 32'b00111111100101111011111101100100, 32'b00111111100101111101010111100100, 32'b00111111100101111110110001101011, 32'b00111111100110000000001011111001, 32'b00111111100110000001100110001101, 32'b00111111100110000011000000101000, 32'b00111111100110000100011011001010, 32'b00111111100110000101110101110010, 32'b00111111100110000111010000100001, 32'b00111111100110001000101011010111, 32'b00111111100110001010000110010100, 32'b00111111100110001011100001010111, 32'b00111111100110001100111100100001, 32'b00111111100110001110010111110010, 32'b00111111100110001111110011001010, 32'b00111111100110010001001110101001, 32'b00111111100110010010101010001111, 32'b00111111100110010100000101111011, 32'b00111111100110010101100001101110, 32'b00111111100110010110111101101000, 32'b00111111100110011000011001101001, 32'b00111111100110011001110101110001, 32'b00111111100110011011010010000000, 32'b00111111100110011100101110010110, 32'b00111111100110011110001010110011, 32'b00111111100110011111100111010110, 32'b00111111100110100001000100000001, 32'b00111111100110100010100000110011, 32'b00111111100110100011111101101011, 32'b00111111100110100101011010101011, 32'b00111111100110100110110111110001, 32'b00111111100110101000010100111111, 32'b00111111100110101001110010010100, 32'b00111111100110101011001111101111, 32'b00111111100110101100101101010010, 32'b00111111100110101110001010111100, 32'b00111111100110101111101000101101, 32'b00111111100110110001000110100101, 32'b00111111100110110010100100100100, 32'b00111111100110110100000010101010, 32'b00111111100110110101100000111000, 32'b00111111100110110110111111001100, 32'b00111111100110111000011101101000, 32'b00111111100110111001111100001011, 32'b00111111100110111011011010110101, 32'b00111111100110111100111001100110, 32'b00111111100110111110011000011111, 32'b00111111100110111111110111011111, 32'b00111111100111000001010110100110, 32'b00111111100111000010110101110100, 32'b00111111100111000100010101001001, 32'b00111111100111000101110100100110, 32'b00111111100111000111010100001010, 32'b00111111100111001000110011110110, 32'b00111111100111001010010011101000, 32'b00111111100111001011110011100010, 32'b00111111100111001101010011100100, 32'b00111111100111001110110011101100, 32'b00111111100111010000010011111100, 32'b00111111100111010001110100010100, 32'b00111111100111010011010100110011, 32'b00111111100111010100110101011001, 32'b00111111100111010110010110000111, 32'b00111111100111010111110110111100, 32'b00111111100111011001010111111001, 32'b00111111100111011010111000111101, 32'b00111111100111011100011010001000, 32'b00111111100111011101111011011011, 32'b00111111100111011111011100110110, 32'b00111111100111100000111110011000, 32'b00111111100111100010100000000001, 32'b00111111100111100100000001110010, 32'b00111111100111100101100011101011, 32'b00111111100111100111000101101011, 32'b00111111100111101000100111110011, 32'b00111111100111101010001010000011, 32'b00111111100111101011101100011010, 32'b00111111100111101101001110111000, 32'b00111111100111101110110001011111, 32'b00111111100111110000010100001101, 32'b00111111100111110001110111000010, 32'b00111111100111110011011010000000, 32'b00111111100111110100111101000101, 32'b00111111100111110110100000010010, 32'b00111111100111111000000011100110, 32'b00111111100111111001100111000010, 32'b00111111100111111011001010100110, 32'b00111111100111111100101110010010, 32'b00111111100111111110010010000101, 32'b00111111100111111111110110000001, 32'b00111111101000000001011010000100, 32'b00111111101000000010111110001111, 32'b00111111101000000100100010100010, 32'b00111111101000000110000110111100, 32'b00111111101000000111101011011111, 32'b00111111101000001001010000001001, 32'b00111111101000001010110100111100, 32'b00111111101000001100011001110110, 32'b00111111101000001101111110111000, 32'b00111111101000001111100100000010, 32'b00111111101000010001001001010100, 32'b00111111101000010010101110101110, 32'b00111111101000010100010100010000, 32'b00111111101000010101111001111010, 32'b00111111101000010111011111101100, 32'b00111111101000011001000101100110, 32'b00111111101000011010101011101000, 32'b00111111101000011100010001110010, 32'b00111111101000011101111000000100, 32'b00111111101000011111011110011111, 32'b00111111101000100001000101000001, 32'b00111111101000100010101011101100, 32'b00111111101000100100010010011110, 32'b00111111101000100101111001011001, 32'b00111111101000100111100000011100, 32'b00111111101000101001000111100111, 32'b00111111101000101010101110111011, 32'b00111111101000101100010110010110, 32'b00111111101000101101111101111010, 32'b00111111101000101111100101100110, 32'b00111111101000110001001101011010, 32'b00111111101000110010110101010111, 32'b00111111101000110100011101011100, 32'b00111111101000110110000101101001, 32'b00111111101000110111101101111110, 32'b00111111101000111001010110011100, 32'b00111111101000111010111111000010, 32'b00111111101000111100100111110001, 32'b00111111101000111110010000101000, 32'b00111111101000111111111001100111, 32'b00111111101001000001100010101111, 32'b00111111101001000011001011111111, 32'b00111111101001000100110101010111, 32'b00111111101001000110011110111000, 32'b00111111101001001000001000100010, 32'b00111111101001001001110010010100, 32'b00111111101001001011011100001110, 32'b00111111101001001101000110010001, 32'b00111111101001001110110000011101, 32'b00111111101001010000011010110001, 32'b00111111101001010010000101001110, 32'b00111111101001010011101111110011, 32'b00111111101001010101011010100001, 32'b00111111101001010111000101010111, 32'b00111111101001011000110000010110, 32'b00111111101001011010011011011110, 32'b00111111101001011100000110101111, 32'b00111111101001011101110010001000, 32'b00111111101001011111011101101010, 32'b00111111101001100001001001010100, 32'b00111111101001100010110101001000, 32'b00111111101001100100100001000100, 32'b00111111101001100110001101001001, 32'b00111111101001100111111001010110, 32'b00111111101001101001100101101101, 32'b00111111101001101011010010001100, 32'b00111111101001101100111110110100, 32'b00111111101001101110101011100101, 32'b00111111101001110000011000011111, 32'b00111111101001110010000101100001, 32'b00111111101001110011110010101101, 32'b00111111101001110101100000000001, 32'b00111111101001110111001101011111, 32'b00111111101001111000111011000101, 32'b00111111101001111010101000110101, 32'b00111111101001111100010110101101, 32'b00111111101001111110000100101111, 32'b00111111101001111111110010111001, 32'b00111111101010000001100001001100, 32'b00111111101010000011001111101001, 32'b00111111101010000100111110001110, 32'b00111111101010000110101100111101, 32'b00111111101010001000011011110101, 32'b00111111101010001010001010110110, 32'b00111111101010001011111010000000, 32'b00111111101010001101101001010011, 32'b00111111101010001111011000110000, 32'b00111111101010010001001000010101, 32'b00111111101010010010111000000100, 32'b00111111101010010100100111111100, 32'b00111111101010010110010111111101, 32'b00111111101010011000001000001000, 32'b00111111101010011001111000011100, 32'b00111111101010011011101000111001, 32'b00111111101010011101011001100000, 32'b00111111101010011111001010001111, 32'b00111111101010100000111011001001, 32'b00111111101010100010101100001011, 32'b00111111101010100100011101010111, 32'b00111111101010100110001110101101, 32'b00111111101010101000000000001100, 32'b00111111101010101001110001110100, 32'b00111111101010101011100011100110, 32'b00111111101010101101010101100001, 32'b00111111101010101111000111100110, 32'b00111111101010110000111001110100, 32'b00111111101010110010101100001100, 32'b00111111101010110100011110101101, 32'b00111111101010110110010001011000, 32'b00111111101010111000000100001101, 32'b00111111101010111001110111001011, 32'b00111111101010111011101010010011, 32'b00111111101010111101011101100101, 32'b00111111101010111111010001000000, 32'b00111111101011000001000100100101, 32'b00111111101011000010111000010011, 32'b00111111101011000100101100001100, 32'b00111111101011000110100000001110, 32'b00111111101011001000010100011010, 32'b00111111101011001010001000101111, 32'b00111111101011001011111101001111, 32'b00111111101011001101110001111000, 32'b00111111101011001111100110101011, 32'b00111111101011010001011011101000, 32'b00111111101011010011010000101111, 32'b00111111101011010101000110000000, 32'b00111111101011010110111011011011, 32'b00111111101011011000110001000000, 32'b00111111101011011010100110101110, 32'b00111111101011011100011100100111, 32'b00111111101011011110010010101010, 32'b00111111101011100000001000110110, 32'b00111111101011100001111111001101, 32'b00111111101011100011110101101110, 32'b00111111101011100101101100011001, 32'b00111111101011100111100011001110, 32'b00111111101011101001011010001101, 32'b00111111101011101011010001010111, 32'b00111111101011101101001000101010, 32'b00111111101011101111000000001000, 32'b00111111101011110000110111110000, 32'b00111111101011110010101111100010, 32'b00111111101011110100100111011110, 32'b00111111101011110110011111100101, 32'b00111111101011111000010111110110, 32'b00111111101011111010010000010001, 32'b00111111101011111100001000110111, 32'b00111111101011111110000001100111, 32'b00111111101011111111111010100001, 32'b00111111101100000001110011100110, 32'b00111111101100000011101100110101, 32'b00111111101100000101100110001110, 32'b00111111101100000111011111110011, 32'b00111111101100001001011001100001, 32'b00111111101100001011010011011010, 32'b00111111101100001101001101011110, 32'b00111111101100001111000111101100, 32'b00111111101100010001000010000100, 32'b00111111101100010010111100101000, 32'b00111111101100010100110111010110, 32'b00111111101100010110110010001110, 32'b00111111101100011000101101010001, 32'b00111111101100011010101000011111, 32'b00111111101100011100100011111000, 32'b00111111101100011110011111011011, 32'b00111111101100100000011011001001, 32'b00111111101100100010010111000010, 32'b00111111101100100100010011000101, 32'b00111111101100100110001111010011, 32'b00111111101100101000001011101101, 32'b00111111101100101010001000010001, 32'b00111111101100101100000100111111, 32'b00111111101100101110000001111001, 32'b00111111101100101111111110111110, 32'b00111111101100110001111100001110, 32'b00111111101100110011111001101000, 32'b00111111101100110101110111001110, 32'b00111111101100110111110100111110, 32'b00111111101100111001110010111010, 32'b00111111101100111011110001000001, 32'b00111111101100111101101111010010, 32'b00111111101100111111101101101111, 32'b00111111101101000001101100010111, 32'b00111111101101000011101011001010, 32'b00111111101101000101101010001000, 32'b00111111101101000111101001010010, 32'b00111111101101001001101000100111, 32'b00111111101101001011101000000111, 32'b00111111101101001101100111110010, 32'b00111111101101001111100111101000, 32'b00111111101101010001100111101010, 32'b00111111101101010011100111110111, 32'b00111111101101010101101000001111, 32'b00111111101101010111101000110011, 32'b00111111101101011001101001100010, 32'b00111111101101011011101010011101, 32'b00111111101101011101101011100011, 32'b00111111101101011111101100110101, 32'b00111111101101100001101110010010, 32'b00111111101101100011101111111010, 32'b00111111101101100101110001101110, 32'b00111111101101100111110011101110, 32'b00111111101101101001110101111001, 32'b00111111101101101011111000010000, 32'b00111111101101101101111010110011, 32'b00111111101101101111111101100001, 32'b00111111101101110010000000011011, 32'b00111111101101110100000011100000, 32'b00111111101101110110000110110010, 32'b00111111101101111000001010001111, 32'b00111111101101111010001101111000, 32'b00111111101101111100010001101100, 32'b00111111101101111110010101101101, 32'b00111111101110000000011001111001, 32'b00111111101110000010011110010010, 32'b00111111101110000100100010110110, 32'b00111111101110000110100111100110, 32'b00111111101110001000101100100010, 32'b00111111101110001010110001101010, 32'b00111111101110001100110110111110, 32'b00111111101110001110111100011110, 32'b00111111101110010001000010001010, 32'b00111111101110010011001000000011, 32'b00111111101110010101001110000111, 32'b00111111101110010111010100011000, 32'b00111111101110011001011010110100, 32'b00111111101110011011100001011101, 32'b00111111101110011101101000010010, 32'b00111111101110011111101111010100, 32'b00111111101110100001110110100001, 32'b00111111101110100011111101111011, 32'b00111111101110100110000101100010, 32'b00111111101110101000001101010100, 32'b00111111101110101010010101010011, 32'b00111111101110101100011101011110, 32'b00111111101110101110100101110110, 32'b00111111101110110000101110011011, 32'b00111111101110110010110111001011, 32'b00111111101110110101000000001000, 32'b00111111101110110111001001010010, 32'b00111111101110111001010010101001, 32'b00111111101110111011011100001100, 32'b00111111101110111101100101111011, 32'b00111111101110111111101111110111, 32'b00111111101111000001111010000000, 32'b00111111101111000100000100010110, 32'b00111111101111000110001110111000, 32'b00111111101111001000011001100111, 32'b00111111101111001010100100100011, 32'b00111111101111001100101111101011, 32'b00111111101111001110111011000001, 32'b00111111101111010001000110100011, 32'b00111111101111010011010010010010, 32'b00111111101111010101011110001111, 32'b00111111101111010111101010011000, 32'b00111111101111011001110110101110, 32'b00111111101111011100000011010001, 32'b00111111101111011110010000000001, 32'b00111111101111100000011100111110, 32'b00111111101111100010101010001000, 32'b00111111101111100100110111100000, 32'b00111111101111100111000101000100, 32'b00111111101111101001010010110110, 32'b00111111101111101011100000110101, 32'b00111111101111101101101111000001, 32'b00111111101111101111111101011010, 32'b00111111101111110010001100000001, 32'b00111111101111110100011010110101, 32'b00111111101111110110101001110110, 32'b00111111101111111000111001000101, 32'b00111111101111111011001000100001, 32'b00111111101111111101011000001010, 32'b00111111101111111111101000000001, 32'b00111111110000000001111000000110, 32'b00111111110000000100001000011000, 32'b00111111110000000110011000111000, 32'b00111111110000001000101001100101, 32'b00111111110000001010111010100000, 32'b00111111110000001101001011101000, 32'b00111111110000001111011100111110, 32'b00111111110000010001101110100010, 32'b00111111110000010100000000010011, 32'b00111111110000010110010010010011, 32'b00111111110000011000100100100000, 32'b00111111110000011010110110111011, 32'b00111111110000011101001001100100, 32'b00111111110000011111011100011010, 32'b00111111110000100001101111011111, 32'b00111111110000100100000010110001, 32'b00111111110000100110010110010010, 32'b00111111110000101000101010000000, 32'b00111111110000101010111101111101, 32'b00111111110000101101010010001000, 32'b00111111110000101111100110100000, 32'b00111111110000110001111011000111, 32'b00111111110000110100001111111100, 32'b00111111110000110110100101000000, 32'b00111111110000111000111010010001, 32'b00111111110000111011001111110001, 32'b00111111110000111101100101011111, 32'b00111111110000111111111011011011, 32'b00111111110001000010010001100110, 32'b00111111110001000100100111111111, 32'b00111111110001000110111110100111, 32'b00111111110001001001010101011101, 32'b00111111110001001011101100100001, 32'b00111111110001001110000011110100, 32'b00111111110001010000011011010110, 32'b00111111110001010010110011000110, 32'b00111111110001010101001011000101, 32'b00111111110001010111100011010010, 32'b00111111110001011001111011101111, 32'b00111111110001011100010100011001, 32'b00111111110001011110101101010011, 32'b00111111110001100001000110011011, 32'b00111111110001100011011111110011, 32'b00111111110001100101111001011001, 32'b00111111110001101000010011001110, 32'b00111111110001101010101101010010, 32'b00111111110001101101000111100100, 32'b00111111110001101111100010000110, 32'b00111111110001110001111100110111, 32'b00111111110001110100010111110111, 32'b00111111110001110110110011000110, 32'b00111111110001111001001110100100, 32'b00111111110001111011101010010010, 32'b00111111110001111110000110001110, 32'b00111111110010000000100010011010, 32'b00111111110010000010111110110101, 32'b00111111110010000101011011011111, 32'b00111111110010000111111000011001, 32'b00111111110010001010010101100010, 32'b00111111110010001100110010111010, 32'b00111111110010001111010000100010, 32'b00111111110010010001101110011001, 32'b00111111110010010100001100100000, 32'b00111111110010010110101010110111, 32'b00111111110010011001001001011101, 32'b00111111110010011011101000010010, 32'b00111111110010011110000111010111, 32'b00111111110010100000100110101100, 32'b00111111110010100011000110010001, 32'b00111111110010100101100110000110, 32'b00111111110010101000000110001010, 32'b00111111110010101010100110011110, 32'b00111111110010101101000111000010, 32'b00111111110010101111100111110110, 32'b00111111110010110010001000111010, 32'b00111111110010110100101010001101, 32'b00111111110010110111001011110001, 32'b00111111110010111001101101100101, 32'b00111111110010111100001111101001, 32'b00111111110010111110110001111101, 32'b00111111110011000001010100100010, 32'b00111111110011000011110111010110, 32'b00111111110011000110011010011011, 32'b00111111110011001000111101110000, 32'b00111111110011001011100001010110, 32'b00111111110011001110000101001011, 32'b00111111110011010000101001010001, 32'b00111111110011010011001101101000, 32'b00111111110011010101110010001111, 32'b00111111110011011000010111000111, 32'b00111111110011011010111100001111, 32'b00111111110011011101100001101000, 32'b00111111110011100000000111010001, 32'b00111111110011100010101101001011, 32'b00111111110011100101010011010110, 32'b00111111110011100111111001110001, 32'b00111111110011101010100000011110, 32'b00111111110011101101000111011011, 32'b00111111110011101111101110101001, 32'b00111111110011110010010110001000, 32'b00111111110011110100111101111000, 32'b00111111110011110111100101111001, 32'b00111111110011111010001110001011, 32'b00111111110011111100110110101110, 32'b00111111110011111111011111100010, 32'b00111111110100000010001000100111, 32'b00111111110100000100110001111110, 32'b00111111110100000111011011100101, 32'b00111111110100001010000101011110, 32'b00111111110100001100101111101001, 32'b00111111110100001111011010000100, 32'b00111111110100010010000100110010, 32'b00111111110100010100101111110000, 32'b00111111110100010111011011000000, 32'b00111111110100011010000110100010, 32'b00111111110100011100110010010101, 32'b00111111110100011111011110011001, 32'b00111111110100100010001010110000, 32'b00111111110100100100110111011000, 32'b00111111110100100111100100010010, 32'b00111111110100101010010001011101, 32'b00111111110100101100111110111011, 32'b00111111110100101111101100101010, 32'b00111111110100110010011010101011, 32'b00111111110100110101001000111111, 32'b00111111110100110111110111100100, 32'b00111111110100111010100110011011, 32'b00111111110100111101010101100100, 32'b00111111110101000000000101000000, 32'b00111111110101000010110100101101, 32'b00111111110101000101100100101101, 32'b00111111110101001000010100111111, 32'b00111111110101001011000101100100, 32'b00111111110101001101110110011010, 32'b00111111110101010000100111100100, 32'b00111111110101010011011000111111, 32'b00111111110101010110001010101101, 32'b00111111110101011000111100101110, 32'b00111111110101011011101111000001, 32'b00111111110101011110100001100111, 32'b00111111110101100001010100011111, 32'b00111111110101100100000111101011, 32'b00111111110101100110111011001000, 32'b00111111110101101001101110111001, 32'b00111111110101101100100010111101, 32'b00111111110101101111010111010011, 32'b00111111110101110010001011111101, 32'b00111111110101110101000000111001, 32'b00111111110101110111110110001001, 32'b00111111110101111010101011101011, 32'b00111111110101111101100001100001, 32'b00111111110110000000010111101010, 32'b00111111110110000011001110000110, 32'b00111111110110000110000100110101, 32'b00111111110110001000111011111000, 32'b00111111110110001011110011001110, 32'b00111111110110001110101010111000, 32'b00111111110110010001100010110101, 32'b00111111110110010100011011000101, 32'b00111111110110010111010011101001, 32'b00111111110110011010001100100001, 32'b00111111110110011101000101101100, 32'b00111111110110011111111111001011, 32'b00111111110110100010111000111110, 32'b00111111110110100101110011000101, 32'b00111111110110101000101101011111, 32'b00111111110110101011101000001110, 32'b00111111110110101110100011010000, 32'b00111111110110110001011110100110, 32'b00111111110110110100011010010001, 32'b00111111110110110111010110001111, 32'b00111111110110111010010010100010, 32'b00111111110110111101001111001001, 32'b00111111110111000000001100000100, 32'b00111111110111000011001001010011, 32'b00111111110111000110000110110111, 32'b00111111110111001001000100101111, 32'b00111111110111001100000010111100, 32'b00111111110111001111000001011101, 32'b00111111110111010010000000010011, 32'b00111111110111010100111111011110, 32'b00111111110111010111111110111101, 32'b00111111110111011010111110110001, 32'b00111111110111011101111110111001, 32'b00111111110111100000111111010111, 32'b00111111110111100100000000001001, 32'b00111111110111100111000001010000, 32'b00111111110111101010000010101100, 32'b00111111110111101101000100011110, 32'b00111111110111110000000110100100, 32'b00111111110111110011001001000000, 32'b00111111110111110110001011110000, 32'b00111111110111111001001110110110, 32'b00111111110111111100010010010010, 32'b00111111110111111111010110000011, 32'b00111111111000000010011010001001, 32'b00111111111000000101011110100100, 32'b00111111111000001000100011010101, 32'b00111111111000001011101000011100, 32'b00111111111000001110101101111001, 32'b00111111111000010001110011101011, 32'b00111111111000010100111001110010, 32'b00111111111000011000000000010000, 32'b00111111111000011011000111000100, 32'b00111111111000011110001110001101, 32'b00111111111000100001010101101101, 32'b00111111111000100100011101100010, 32'b00111111111000100111100101101110, 32'b00111111111000101010101110001111, 32'b00111111111000101101110111000111, 32'b00111111111000110001000000010110, 32'b00111111111000110100001001111010, 32'b00111111111000110111010011110101, 32'b00111111111000111010011110000111, 32'b00111111111000111101101000101110, 32'b00111111111001000000110011101101, 32'b00111111111001000011111111000010, 32'b00111111111001000111001010101110, 32'b00111111111001001010010110110000, 32'b00111111111001001101100011001001, 32'b00111111111001010000101111111010, 32'b00111111111001010011111101000001, 32'b00111111111001010111001010011111, 32'b00111111111001011010011000010100, 32'b00111111111001011101100110100000, 32'b00111111111001100000110101000011, 32'b00111111111001100100000011111110, 32'b00111111111001100111010011010000, 32'b00111111111001101010100010111001, 32'b00111111111001101101110010111010, 32'b00111111111001110001000011010010, 32'b00111111111001110100010100000001, 32'b00111111111001110111100101001001, 32'b00111111111001111010110110100111, 32'b00111111111001111110001000011110, 32'b00111111111010000001011010101100, 32'b00111111111010000100101101010011, 32'b00111111111010001000000000010001, 32'b00111111111010001011010011100111, 32'b00111111111010001110100111010101, 32'b00111111111010010001111011011011, 32'b00111111111010010101001111111010, 32'b00111111111010011000100100110000, 32'b00111111111010011011111001111111, 32'b00111111111010011111001111100110, 32'b00111111111010100010100101100110, 32'b00111111111010100101111011111110, 32'b00111111111010101001010010101111, 32'b00111111111010101100101001111000, 32'b00111111111010110000000001011010, 32'b00111111111010110011011001010101, 32'b00111111111010110110110001101001, 32'b00111111111010111010001010010101, 32'b00111111111010111101100011011011, 32'b00111111111011000000111100111001, 32'b00111111111011000100010110110001, 32'b00111111111011000111110001000010, 32'b00111111111011001011001011101100, 32'b00111111111011001110100110101111, 32'b00111111111011010010000010001011, 32'b00111111111011010101011110000010, 32'b00111111111011011000111010010001, 32'b00111111111011011100010110111010, 32'b00111111111011011111110011111101, 32'b00111111111011100011010001011001, 32'b00111111111011100110101111010000, 32'b00111111111011101010001101100000, 32'b00111111111011101101101100001010, 32'b00111111111011110001001011001110, 32'b00111111111011110100101010101100, 32'b00111111111011111000001010100100, 32'b00111111111011111011101010110110, 32'b00111111111011111111001011100011, 32'b00111111111100000010101100101010, 32'b00111111111100000110001110001100, 32'b00111111111100001001110000001000, 32'b00111111111100001101010010011110, 32'b00111111111100010000110101001111, 32'b00111111111100010100011000011011, 32'b00111111111100010111111100000010, 32'b00111111111100011011100000000011, 32'b00111111111100011111000100100000, 32'b00111111111100100010101001010111, 32'b00111111111100100110001110101010, 32'b00111111111100101001110100011000, 32'b00111111111100101101011010100001, 32'b00111111111100110001000001000101, 32'b00111111111100110100101000000101, 32'b00111111111100111000001111100000, 32'b00111111111100111011110111010111, 32'b00111111111100111111011111101001, 32'b00111111111101000011001000010111, 32'b00111111111101000110110001100001, 32'b00111111111101001010011011000110, 32'b00111111111101001110000101001000, 32'b00111111111101010001101111100101, 32'b00111111111101010101011010011111, 32'b00111111111101011001000101110101, 32'b00111111111101011100110001100111, 32'b00111111111101100000011101110101, 32'b00111111111101100100001010100000, 32'b00111111111101100111110111100111, 32'b00111111111101101011100101001011, 32'b00111111111101101111010011001100, 32'b00111111111101110011000001101001, 32'b00111111111101110110110000100011, 32'b00111111111101111010011111111010, 32'b00111111111101111110001111101110, 32'b00111111111110000001111111111111, 32'b00111111111110000101110000101101, 32'b00111111111110001001100001111000, 32'b00111111111110001101010011100001, 32'b00111111111110010001000101100111, 32'b00111111111110010100111000001010, 32'b00111111111110011000101011001011, 32'b00111111111110011100011110101010, 32'b00111111111110100000010010100110, 32'b00111111111110100100000111000001, 32'b00111111111110100111111011111001, 32'b00111111111110101011110001001111, 32'b00111111111110101111100111000011, 32'b00111111111110110011011101010101, 32'b00111111111110110111010100000110, 32'b00111111111110111011001011010101, 32'b00111111111110111111000011000010, 32'b00111111111111000010111011001110, 32'b00111111111111000110110011111000, 32'b00111111111111001010101101000001, 32'b00111111111111001110100110101001, 32'b00111111111111010010100000101111, 32'b00111111111111010110011011010101, 32'b00111111111111011010010110011010, 32'b00111111111111011110010001111101, 32'b00111111111111100010001110000000, 32'b00111111111111100110001010100011, 32'b00111111111111101010000111100100, 32'b00111111111111101110000101000110, 32'b00111111111111110010000011000110, 32'b00111111111111110110000001100111, 32'b00111111111111111010000000100111, 32'b00111111111111111110000000000111};

    wire [9:0] key0;
    assign key0 = x[22:13];
    wire [31:0] ax2; 
    wire [31:0] test_a0;
    wire [31:0] test_b0;

    assign test_a0 = a_table[key0];
    assign test_b0 = b_table[key0];
    wire [31:0] x_m0;
    assign x_m0 = {1'b0, 8'd127, x[22:0]};
    fmul fmull(test_a0,x_m0,ax2,clk);
    reg [31:0] ax_3;
    reg[31:0] x_1;
    reg[31:0] x_2;
    reg[31:0] x_3;
    reg[31:0] x_4;
    reg[31:0] x_5;


    reg [31:0] test_b_1;
    reg [31:0] test_b_2;
    reg [31:0] test_b_3;
    
    always @(posedge clk) begin
      ax_3<=ax2;
      x_1<=x;
      x_2<=x_1;
      x_3<=x_2;
      x_4<=x_3;
      x_5<=x_4;

      test_b_1<=test_b0;
      test_b_2<=test_b_1;
      test_b_3<=test_b_2;

   end
    wire [31:0] y_sub5;
    fadd faddd(test_b_3,ax_3,y_sub5,clk);
    wire [31:0] y_sub55;
    wire [7:0] y_sub_e;
    assign y_sub_e =  y_sub5[30:23] - (x_5[30:23] - 8'd127);
    assign y_sub55 = {x_5[31:31],y_sub_e, y_sub5[22:0] };
    assign y = (x_5[30:23]==0) ? 32'b01111111100000000000000000000000 : y_sub55;
endmodule

module fdiv (input wire [31:0] x1,
             input wire [31:0] x2,
             output wire [31:0] y,
              input wire clk);

   reg [31:0] x1_1;
   reg [31:0] x2_1;

   always @(posedge clk) begin
      x1_1<=x1;
      x2_1<=x2;
   end
    
    wire [31:0] x_m1_1;
    reg [31:0] x_m1_2;
    reg [31:0] x_m1_3;
    reg [31:0] x_m1_4;
    reg [31:0] x_m1_5;
    reg [31:0] x_m1_6;


    assign x_m1_1 = {1'b0, 8'd127, x1_1[22:0]};
    wire [31:0] x_m2_1;
    assign x_m2_1 = {1'b0, 8'd127, x2_1[22:0]};
    wire [31:0] inv_x_m2_6;
    finv finvv(x_m2_1, inv_x_m2_6,clk);
    wire [31:0] m1m2_8;
    always @(posedge clk) begin
      x_m1_2<=x_m1_1;
      x_m1_3<=x_m1_2;
      x_m1_4<=x_m1_3;
      x_m1_5<=x_m1_4;
      x_m1_6<=x_m1_5;
   end
   reg [31:0] x1_2;
   reg [31:0] x2_2;
   reg [31:0] x1_3;
   reg [31:0] x2_3;
   reg [31:0] x1_4;
   reg [31:0] x2_4;
   reg [31:0] x1_5;
   reg [31:0] x2_5;
   reg [31:0] x1_6;
   reg [31:0] x2_6;
   reg [31:0] x1_7;
   reg [31:0] x2_7;
   reg [31:0] x1_8;
   reg [31:0] x2_8;
  
    fmul fmull(x_m1_6,inv_x_m2_6,m1m2_8,clk);
    always @(posedge clk) begin
       x1_2<=x1_1;
       x2_2<=x2_1;
       x1_3<=x1_2;
       x2_3<=x2_2;
       x1_4<=x1_3;
       x2_4<=x2_3;
       x1_5<=x1_4;
       x2_5<=x2_4;
       x1_6<=x1_5;
       x2_6<=x2_5;
       x1_7<=x1_6;
       x2_7<=x2_6;
       x1_8<=x1_7;
       x2_8<=x2_7;

   end
    wire [7:0] ey;
    assign ey = (m1m2_8[30:23]==127) ? x1_8[30:23]-x2_8[30:23] +127: x1_8[30:23]-x2_8[30:23]+126;
    wire sy;
    assign sy = x1_8[31:31] ^ x2_8[31:31];
    wire [31:0] y_sub;
    assign y_sub = {sy, ey, m1m2_8[22:0]};
    assign y = (x1_8[30:23]==0) ? 32'b0 : (x2_8[30:23]==0) ? 32'b01111111100000000000000000000000 : y_sub;


endmodule